* NGSPICE file created from asic_flat.ext - technology: sky130A

.subckt asic_flat ua[0] ua[1] ua[2] ua[3] ua[4] ua[5] VGND VAPWR
X0 a_9577_9007.t4 a_9039_8199.t2 a_9039_8199.t3 VAPWR.t28 sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=2.5 l=2.4
**devattr s=29000,1116 d=29000,1116
X1 VGND.t78 VGND.t86 BIAS_1_0.XQ12.Emitter sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X2 a_3378_41806# a_3378_35748# VGND.t7 sky130_fd_pr__res_xhigh_po_0p35 l=25
X3 VAPWR.t8 ua[5].t0 a_12179_10665# VAPWR.t7 sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.145 ps=1.29 w=1 l=0.5
**devattr s=5800,258 d=5800,258
X4 a_4562_41806# a_4858_35748# VGND.t31 sky130_fd_pr__res_xhigh_po_0p35 l=25
X5 a_2786_41806# a_2786_35748# VGND.t21 sky130_fd_pr__res_xhigh_po_0p35 l=25
X6 a_5450_35748# a_5450_30348# VGND.t10 sky130_fd_pr__res_xhigh_po_0p35 l=25
X7 Timming_0.Vd.t23 a_16597_7688.t14 a_16597_7688.t15 VGND.t104 sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=10 l=0.5
**devattr s=58000,2058 d=58000,2058
X8 VCR_0.VT.t9 ua[2].t2 VGND.t56 VGND.t55 sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=5 l=1
**devattr s=29000,1058 d=29000,1058
X9 a_7586_26267# a_9886_26267# VGND.t6 sky130_fd_pr__res_xhigh_po_0p35 l=9.5
X10 a_9886_25971# a_12844_25971# VGND.t1 sky130_fd_pr__res_xhigh_po_0p35 l=9.5
X11 a_10404_14647.t6 a_6404_16954.t4 a_6404_16954.t5 VAPWR.t1 sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=10 l=20
**devattr s=116000,4116 d=116000,4116
X12 VGND.t24 ua[2].t3 VCR_0.VT.t8 VGND.t23 sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=5 l=1
**devattr s=29000,1058 d=29000,1058
X13 Timming_0.Vd.t22 a_16597_7688.t20 a_16597_7688.t21 VGND.t54 sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=10 l=0.5
**devattr s=58000,2058 d=58000,2058
X14 a_12495_10665# latch_sch_0.Qn.t4 VAPWR.t37 VAPWR.t36 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=0.5
**devattr s=5800,258 d=5800,258
X15 ua[0].t7 a_21737_7899.t3 VAPWR.t10 VAPWR.t9 sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=8.5 l=1
**devattr s=49300,1758 d=49300,1758
X16 a_7586_27451# a_9886_27747# VGND.t6 sky130_fd_pr__res_xhigh_po_0p35 l=9.5
X17 VGND.t73 a_5453_6051.t3 a_5453_6051.t4 VGND.t35 sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=6
**devattr s=11600,516 d=11600,516
X18 a_5154_35748# a_4858_30348# VGND.t72 sky130_fd_pr__res_xhigh_po_0p35 l=25
X19 ua[0].t6 a_21737_7899.t4 VAPWR.t17 VAPWR.t16 sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=8.5 l=1
**devattr s=98600,3516 d=49300,1758
X20 a_3082_35748# a_3082_30348# VGND.t9 sky130_fd_pr__res_xhigh_po_0p35 l=25
X21 a_4562_35748# a_4266_30348# VGND.t17 sky130_fd_pr__res_xhigh_po_0p35 l=25
X22 latch_sch_0.R.t0 a_5453_6051.t8 VGND.t43 VGND.t42 sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=2.2
**devattr s=11600,516 d=11600,516
X23 a_3970_35748# a_3674_30348# VGND.t16 sky130_fd_pr__res_xhigh_po_0p35 l=25
X24 a_9886_27451# a_12844_27155# VGND.t1 sky130_fd_pr__res_xhigh_po_0p35 l=9.5
X25 VGND.t78 VGND.t85 BIAS_1_0.XQ12.Emitter sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X26 a_6404_16954.t3 a_6404_16954.t2 a_10404_14647.t5 VAPWR.t3 sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=10 l=20
**devattr s=116000,4116 d=116000,4116
X27 a_7586_25083# a_9886_25379# VGND.t6 sky130_fd_pr__res_xhigh_po_0p35 l=9.5
X28 VGND.t67 a_5453_6051.t9 a_5453_6767.t3 VGND.t35 sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=6
**devattr s=11600,516 d=11600,516
X29 VGND.t78 VGND.t84 BIAS_1_0.XQ12.Emitter sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X30 a_7586_26859# a_9886_26859# VGND.t6 sky130_fd_pr__res_xhigh_po_0p35 l=9.5
X31 a_20802_14722.t1 VGND.t109 sky130_fd_pr__cap_mim_m3_1 l=27.5 w=27.5
X32 VGND.t78 VGND.t83 BIAS_1_0.XQ12.Emitter sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X33 a_16169_6107# a_15873_2607# VGND.t11 sky130_fd_pr__res_xhigh_po_0p35 l=15.5
X34 a_4266_35748# a_4266_30348# VGND.t8 sky130_fd_pr__res_xhigh_po_0p35 l=25
X35 a_9886_25083# a_11336_20947# VGND.t1 sky130_fd_pr__res_xhigh_po_0p35 l=9.5
X36 a_16597_7688.t39 a_16597_7688.t38 Timming_0.Vd.t21 VGND.t103 sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=10 l=0.5
**devattr s=58000,2058 d=58000,2058
X37 Timming_0.Vd.t20 a_16597_7688.t36 a_16597_7688.t37 VGND.t74 sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=10 l=0.5
**devattr s=58000,2058 d=58000,2058
X38 a_3674_35748# a_3674_30348# VGND.t12 sky130_fd_pr__res_xhigh_po_0p35 l=25
X39 VAPWR.t23 a_21737_7899.t5 ua[0].t5 VAPWR.t22 sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=8.5 l=1
**devattr s=49300,1758 d=49300,1758
X40 a_15873_10265# Timming_0.Vd.t0 VGND.t11 sky130_fd_pr__res_xhigh_po_0p35 l=15.5
X41 a_14097_6107# a_14097_2607# VGND.t106 sky130_fd_pr__res_xhigh_po_0p35 l=15.5
X42 a_5453_6051.t7 COMP_2_0.vin_n.t2 a_6061_11160.t1 VAPWR.t15 sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=2.5 l=2.4
**devattr s=29000,1116 d=29000,1116
X43 a_9886_26563# a_12844_26563# VGND.t1 sky130_fd_pr__res_xhigh_po_0p35 l=9.5
X44 a_14097_10265# a_14097_6107# VGND.t106 sky130_fd_pr__res_xhigh_po_0p35 l=15.5
X45 latch_sch_0.Qn.t3 ua[5].t1 VGND.t64 VGND.t63 sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
**devattr s=11600,516 d=11600,516
X46 a_10404_14647.t0 delay_1_0.vd_n.t1 VAPWR.t5 VAPWR.t4 sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=9.95
**devattr s=11600,516 d=11600,516
X47 VGND.t116 ua[2].t4 VCR_0.VT.t7 VGND.t115 sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=5 l=1
**devattr s=29000,1058 d=29000,1058
X48 a_17267_7131# ua[3].t0 a_17853_5073# VGND.t98 sky130_fd_pr__nfet_05v0_nvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=10
**devattr s=11600,516 d=11600,516
X49 VGND.t129 latch_sch_0.Qn.t5 Timming_0.Vd.t25 VGND.t128 sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
**devattr s=11600,516 d=11600,516
X50 a_19306_5807# a_17853_5073# VGND.t20 sky130_fd_pr__res_xhigh_po_0p35 l=14
X51 a_3378_35748# a_3082_30348# VGND.t7 sky130_fd_pr__res_xhigh_po_0p35 l=25
X52 a_16597_7688.t35 a_16597_7688.t34 Timming_0.Vd.t19 VGND.t48 sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=10 l=0.5
**devattr s=58000,2058 d=58000,2058
X53 a_2786_35748# latch_sch_0.Qn.t0 VGND.t21 sky130_fd_pr__res_xhigh_po_0p35 l=25
X54 a_4858_35748# a_4858_30348# VGND.t31 sky130_fd_pr__res_xhigh_po_0p35 l=25
X55 latch_sch_0.R.t2 a_9039_8199.t5 a_9577_9007.t5 VAPWR.t27 sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=2.5 l=2.4
**devattr s=29000,1116 d=29000,1116
X56 VGND.t18 VGND.t19 VGND.t1 sky130_fd_pr__res_xhigh_po_0p35 l=9.5
X57 a_18714_5807# ua[2].t1 VGND.t130 sky130_fd_pr__res_xhigh_po_0p35 l=14
X58 a_6404_16954.t0 a_11329_22619.t7 a_11336_20947# VGND.t22 sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=1.45 ps=10.58 w=5 l=20
**devattr s=58000,2116 d=58000,2116
X59 a_9886_25675# a_12844_25379# VGND.t1 sky130_fd_pr__res_xhigh_po_0p35 l=9.5
X60 ua[0].t4 a_21737_7899.t6 VAPWR.t21 VAPWR.t20 sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=8.5 l=1
**devattr s=49300,1758 d=49300,1758
X61 a_5453_6767.t7 a_5453_6767.t6 VGND.t75 VGND.t46 sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=6
**devattr s=11600,516 d=11600,516
X62 a_16597_7688.t3 a_16597_7688.t2 Timming_0.Vd.t18 VGND.t114 sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=10 l=0.5
**devattr s=58000,2058 d=58000,2058
X63 Timming_0.Vd.t1 latch_sch_0.R.t3 VGND.t27 VGND.t26 sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
**devattr s=11600,516 d=11600,516
X64 a_17267_7131# ua[3].t1 a_16681_5073# VGND.t51 sky130_fd_pr__nfet_05v0_nvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=10
**devattr s=11600,516 d=11600,516
X65 VGND.t4 Timming_0.Vd.t26 latch_sch_0.Qn.t2 VGND.t3 sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
**devattr s=11600,516 d=11600,516
X66 VGND.t78 VGND.t82 BIAS_1_0.XQ12.Emitter sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X67 a_9886_27155# a_12844_27155# VGND.t1 sky130_fd_pr__res_xhigh_po_0p35 l=9.5
X68 a_11329_22619.t0 a_20802_14722.t2 a_10404_14647.t1 VAPWR.t14 sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=20
**devattr s=5800,316 d=5800,316
X69 a_16597_7688.t41 a_16597_7688.t40 Timming_0.Vd.t17 VGND.t91 sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=10 l=0.5
**devattr s=58000,2058 d=116000,4116
X70 Timming_0.Vd.t16 a_16597_7688.t18 a_16597_7688.t19 VGND.t37 sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=10 l=0.5
**devattr s=58000,2058 d=58000,2058
X71 VGND.t121 VGND.t122 VGND.t1 sky130_fd_pr__res_xhigh_po_0p35 l=9.5
X72 a_10404_14647.t7 a_6404_16954.t6 a_11329_22619.t2 VAPWR.t1 sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=10 l=20
**devattr s=116000,4116 d=116000,4116
X73 a_20802_14722.t3 VGND.t93 sky130_fd_pr__cap_mim_m3_1 l=27.5 w=27.5
X74 VAPWR.t39 a_21737_7899.t7 ua[0].t3 VAPWR.t38 sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=8.5 l=1
**devattr s=49300,1758 d=49300,1758
X75 Timming_0.Vd.t24 latch_sch_0.R.t4 a_12495_10665# VAPWR.t31 sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.145 ps=1.29 w=1 l=0.5
**devattr s=5800,258 d=11600,516
X76 a_16597_7688.t44 ua[3].t2 a_16681_5073# VGND.t76 sky130_fd_pr__nfet_05v0_nvt ad=0 pd=0 as=0.29 ps=2.58 w=1 l=10
**devattr s=11600,516 d=11600,516
X77 a_5453_6051.t5 a_5453_6767.t8 VGND.t47 VGND.t46 sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=6
**devattr s=11600,516 d=11600,516
X78 VGND.t78 VGND.t81 BIAS_1_0.XQ12.Emitter sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X79 delay_1_0.vd_n.t0 VGND.t131 a_8279_30718# VAPWR.t26 sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=10
**devattr s=11600,516 d=11600,516
X80 a_14985_6107# a_15281_2607# VGND.t33 sky130_fd_pr__res_xhigh_po_0p35 l=15.5
X81 a_5453_6767.t0 VCR_0.VT.t11 a_6061_11160.t3 VAPWR.t15 sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=2.5 l=2.4
**devattr s=29000,1116 d=29000,1116
X82 Timming_0.Vd.t15 a_16597_7688.t6 a_16597_7688.t7 VGND.t62 sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=10 l=0.5
**devattr s=58000,2058 d=58000,2058
X83 delay_1_0.vd_n.t2 VGND.t102 sky130_fd_pr__cap_mim_m3_1 l=30 w=30
X84 a_16597_7688.t5 a_16597_7688.t4 Timming_0.Vd.t14 VGND.t59 sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=10 l=0.5
**devattr s=58000,2058 d=58000,2058
X85 Timming_0.Vd.t13 a_16597_7688.t8 a_16597_7688.t9 VGND.t125 sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=10 l=0.5
**devattr s=116000,4116 d=58000,2058
X86 a_15281_10265# a_14985_6765# VGND.t33 sky130_fd_pr__res_xhigh_po_0p35 l=15.5
X87 a_6061_11160.t2 VCR_0.VT.t12 a_5453_6767.t1 VAPWR.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=2.5 l=2.4
**devattr s=29000,1116 d=29000,1116
X88 a_9886_26267# a_12844_25971# VGND.t1 sky130_fd_pr__res_xhigh_po_0p35 l=9.5
X89 VGND.t39 ua[2].t5 VCR_0.VT.t6 VGND.t38 sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=5 l=1
**devattr s=29000,1058 d=58000,2116
X90 a_15577_6107# a_15281_2607# VGND.t32 sky130_fd_pr__res_xhigh_po_0p35 l=15.5
X91 a_14393_6107# a_14097_2607# VGND.t45 sky130_fd_pr__res_xhigh_po_0p35 l=15.5
X92 a_9577_9007.t2 a_9039_8199.t6 latch_sch_0.R.t1 VAPWR.t28 sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=2.5 l=2.4
**devattr s=29000,1116 d=29000,1116
X93 VCR_0.VT.t5 ua[2].t6 VGND.t61 VGND.t60 sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=5 l=1
**devattr s=29000,1058 d=29000,1058
X94 a_15281_10265# a_15577_6765# VGND.t32 sky130_fd_pr__res_xhigh_po_0p35 l=15.5
X95 a_14097_10265# a_14393_6765# VGND.t45 sky130_fd_pr__res_xhigh_po_0p35 l=15.5
X96 a_9886_27747# BIAS_1_0.XQ12.Emitter VGND.t1 sky130_fd_pr__res_xhigh_po_0p35 l=9.5
X97 VGND.t111 ua[2].t7 VCR_0.VT.t4 VGND.t110 sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=5 l=1
**devattr s=29000,1058 d=29000,1058
X98 a_14393_6107# a_14689_2607# VGND.t5 sky130_fd_pr__res_xhigh_po_0p35 l=15.5
X99 a_16597_7688.t17 a_16597_7688.t16 Timming_0.Vd.t12 VGND.t58 sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=10 l=0.5
**devattr s=58000,2058 d=58000,2058
X100 a_8582_24056# COMP_2_0.vb.t4 a_8096_19998# VGND.t30 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=20
**devattr s=5800,316 d=5800,316
X101 a_7586_25675# a_9886_25971# VGND.t6 sky130_fd_pr__res_xhigh_po_0p35 l=9.5
X102 a_7124_24056# COMP_2_0.vb.t5 a_8096_19998# VGND.t49 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=20
**devattr s=5800,316 d=5800,316
X103 VCR_0.VT.t3 ua[2].t8 VGND.t90 VGND.t89 sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=5 l=1
**devattr s=29000,1058 d=29000,1058
X104 ua[0].t2 a_21737_7899.t8 VAPWR.t33 VAPWR.t32 sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=8.5 l=1
**devattr s=49300,1758 d=49300,1758
X105 a_14689_10265# a_14393_6765# VGND.t5 sky130_fd_pr__res_xhigh_po_0p35 l=15.5
X106 VGND.t36 a_5453_6767.t9 a_5453_6051.t0 VGND.t35 sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=6
**devattr s=11600,516 d=11600,516
X107 a_16597_7688.t13 a_16597_7688.t12 Timming_0.Vd.t11 VGND.t97 sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=10 l=0.5
**devattr s=58000,2058 d=58000,2058
X108 Timming_0.Vd.t10 a_16597_7688.t22 a_16597_7688.t23 VGND.t69 sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=10 l=0.5
**devattr s=58000,2058 d=58000,2058
X109 a_9886_25379# a_12844_25379# VGND.t1 sky130_fd_pr__res_xhigh_po_0p35 l=9.5
X110 a_12179_10665# Timming_0.Vd.t27 latch_sch_0.Qn.t1 VAPWR.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=0.5
**devattr s=11600,516 d=5800,258
X111 VGND.t119 a_5453_6767.t10 a_9039_8199.t4 VGND.t118 sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=2.2
**devattr s=11600,516 d=11600,516
X112 a_17267_4669# ua[4].t0 ua[2].t0 VGND.t98 sky130_fd_pr__nfet_05v0_nvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=10
**devattr s=11600,516 d=11600,516
X113 a_9886_26859# a_12844_26563# VGND.t1 sky130_fd_pr__res_xhigh_po_0p35 l=9.5
X114 a_7586_27451# a_9886_27451# VGND.t6 sky130_fd_pr__res_xhigh_po_0p35 l=9.5
X115 a_9554_24056# COMP_2_0.vb.t6 a_9068_19998# VGND.t13 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=20
**devattr s=5800,316 d=5800,316
X116 a_16597_7688.t31 a_16597_7688.t30 Timming_0.Vd.t9 VGND.t34 sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=10 l=0.5
**devattr s=58000,2058 d=58000,2058
X117 a_8582_24056# COMP_2_0.vb.t7 a_9068_19998# VGND.t44 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=20
**devattr s=5800,316 d=5800,316
X118 BIAS_1_0.XQ4.Emitter.t1 a_11329_22619.t3 a_11329_22619.t4 VGND.t22 sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=3 l=20
**devattr s=34800,1316 d=34800,1316
X119 COMP_2_0.vin_n.t1 a_6064_20056# a_6064_20056# VGND.t96 sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.145 ps=1.58 w=0.5 l=20
**devattr s=5800,316 d=5800,316
X120 BIAS_1_0.XQ4.Emitter.t0 a_11329_22619.t5 a_11329_22619.t6 VGND.t107 sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=3 l=20
**devattr s=34800,1316 d=34800,1316
X121 VGND.t113 a_5453_6767.t4 a_5453_6767.t5 VGND.t35 sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=6
**devattr s=11600,516 d=11600,516
X122 a_7586_25083# a_9886_25083# VGND.t6 sky130_fd_pr__res_xhigh_po_0p35 l=9.5
X123 delay_1_0.vd_n.t3 VGND.t0 sky130_fd_pr__cap_mim_m3_1 l=30 w=30
X124 VAPWR.t35 a_21737_7899.t9 ua[0].t1 VAPWR.t34 sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=8.5 l=1
**devattr s=49300,1758 d=49300,1758
X125 a_16597_7688.t1 a_16597_7688.t0 Timming_0.Vd.t8 VGND.t53 sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=10 l=0.5
**devattr s=58000,2058 d=58000,2058
X126 a_16597_7688.t11 a_16597_7688.t10 Timming_0.Vd.t7 VGND.t105 sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=10 l=0.5
**devattr s=58000,2058 d=58000,2058
X127 VGND.t78 VGND.t80 BIAS_1_0.XQ12.Emitter sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X128 a_9554_24056# COMP_2_0.vb.t8 a_10040_19998# VGND.t68 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=20
**devattr s=5800,316 d=5800,316
X129 a_11329_22619.t1 a_6404_16954.t7 a_10404_14647.t3 VAPWR.t3 sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=10 l=20
**devattr s=116000,4116 d=116000,4116
X130 a_20802_14722.t0 VGND.t132 a_10404_14647.t9 VAPWR.t11 sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=20
**devattr s=5800,316 d=5800,316
X131 a_9577_9007.t0 COMP_2_0.vb.t9 a_6061_11160.t4 VAPWR.t13 sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=2 l=20
**devattr s=23200,916 d=23200,916
X132 a_5154_41806# a_5450_35748# VGND.t10 sky130_fd_pr__res_xhigh_po_0p35 l=25
X133 a_7586_26267# a_9886_26563# VGND.t6 sky130_fd_pr__res_xhigh_po_0p35 l=9.5
X134 a_10404_14647.t2 a_6404_16954.t8 COMP_2_0.vb.t1 VAPWR.t6 sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1.5 l=20
**devattr s=17400,716 d=17400,716
X135 a_21737_7899.t0 ua[1].t0 a_21737_5649# VGND.t14 sky130_fd_pr__nfet_05v0_nvt ad=0 pd=0 as=2.9 ps=20.58 w=10 l=9
**devattr s=116000,4116 d=116000,4116
X136 VGND.t41 ua[2].t9 VCR_0.VT.t2 VGND.t40 sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=5 l=1
**devattr s=29000,1058 d=29000,1058
X137 a_17267_4669# ua[4].t1 a_16681_2611# VGND.t51 sky130_fd_pr__nfet_05v0_nvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=10
**devattr s=11600,516 d=11600,516
X138 a_21737_3791# a_21737_7899.t10 VCR_0.VT.t10 VGND.t124 sky130_fd_pr__nfet_05v0_nvt ad=2.9 pd=20.58 as=0 ps=0 w=10 l=9
**devattr s=116000,4116 d=116000,4116
X139 VCR_0.VT.t1 ua[2].t10 VGND.t127 VGND.t126 sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=5 l=1
**devattr s=58000,2116 d=29000,1058
X140 a_7124_24056# COMP_2_0.vb.t2 COMP_2_0.vb.t3 VGND.t120 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=20
**devattr s=5800,316 d=5800,316
X141 a_9039_8199.t1 a_9039_8199.t0 a_9577_9007.t3 VAPWR.t27 sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=2.5 l=2.4
**devattr s=29000,1116 d=29000,1116
X142 a_7124_24056# a_6064_20056# a_6638_19998# VGND.t95 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=20
**devattr s=5800,316 d=5800,316
X143 delay_1_0.vd_n.t4 VGND.t108 sky130_fd_pr__cap_mim_m3_1 l=30 w=30
X144 a_15577_6107# a_15873_2607# VGND.t25 sky130_fd_pr__res_xhigh_po_0p35 l=15.5
X145 a_16169_6107# ua[4].t2 a_16681_2611# VGND.t76 sky130_fd_pr__nfet_05v0_nvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=10
**devattr s=11600,516 d=11600,516
X146 VCR_0.VT.t0 ua[2].t11 VGND.t66 VGND.t65 sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=5 l=1
**devattr s=29000,1058 d=29000,1058
X147 a_2786_41806# a_3082_35748# VGND.t9 sky130_fd_pr__res_xhigh_po_0p35 l=25
X148 a_5154_41806# a_5154_35748# VGND.t72 sky130_fd_pr__res_xhigh_po_0p35 l=25
X149 a_15873_10265# a_15577_6765# VGND.t25 sky130_fd_pr__res_xhigh_po_0p35 l=15.5
X150 a_5453_6767.t2 a_5453_6051.t10 VGND.t92 VGND.t46 sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=6
**devattr s=11600,516 d=11600,516
X151 a_4562_41806# a_4562_35748# VGND.t17 sky130_fd_pr__res_xhigh_po_0p35 l=25
X152 VGND.t70 VGND.t71 VGND.t6 sky130_fd_pr__res_xhigh_po_0p35 l=9.5
X153 a_14985_6107# a_14689_2607# VGND.t15 sky130_fd_pr__res_xhigh_po_0p35 l=15.5
X154 a_3970_41806# a_3970_35748# VGND.t16 sky130_fd_pr__res_xhigh_po_0p35 l=25
X155 a_7586_25675# a_9886_25675# VGND.t6 sky130_fd_pr__res_xhigh_po_0p35 l=9.5
X156 Timming_0.Vd.t6 a_16597_7688.t32 a_16597_7688.t33 VGND.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=10 l=0.5
**devattr s=58000,2058 d=58000,2058
X157 a_21737_7899.t2 a_21737_7899.t1 VAPWR.t30 VAPWR.t29 sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=4 l=1
**devattr s=46400,1716 d=46400,1716
X158 a_14689_10265# a_14985_6765# VGND.t15 sky130_fd_pr__res_xhigh_po_0p35 l=15.5
X159 a_10404_14647.t4 a_6404_16954.t9 COMP_2_0.vb.t0 VAPWR.t6 sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1.5 l=20
**devattr s=17400,716 d=17400,716
X160 Timming_0.Vd.t5 a_16597_7688.t26 a_16597_7688.t27 VGND.t123 sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=10 l=0.5
**devattr s=58000,2058 d=58000,2058
X161 a_16597_7688.t29 a_16597_7688.t28 Timming_0.Vd.t4 VGND.t57 sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=10 l=0.5
**devattr s=58000,2058 d=58000,2058
X162 VGND.t78 VGND.t77 BIAS_1_0.XQ4.Emitter.t2 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X163 a_6404_16954.t1 a_11329_22619.t8 a_11336_20947# VGND.t52 sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=1.45 ps=10.58 w=5 l=20
**devattr s=58000,2116 d=58000,2116
X164 a_9577_9007.t1 delay_1_0.vd_n.t5 VAPWR.t25 VAPWR.t24 sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=10.05
**devattr s=11600,516 d=11600,516
X165 a_3970_41806# a_4266_35748# VGND.t8 sky130_fd_pr__res_xhigh_po_0p35 l=25
X166 delay_1_0.vd_n.t6 VGND.t87 sky130_fd_pr__cap_mim_m3_1 l=30 w=30
X167 a_5453_6051.t2 a_5453_6051.t1 VGND.t117 VGND.t46 sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=6
**devattr s=11600,516 d=11600,516
X168 a_21737_5649# ua[1].t1 a_21737_3791# VGND.t14 sky130_fd_pr__nfet_05v0_nvt ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=9
**devattr s=116000,4116 d=116000,4116
X169 a_3378_41806# a_3674_35748# VGND.t12 sky130_fd_pr__res_xhigh_po_0p35 l=25
X170 COMP_2_0.vin_n.t0 a_6064_20056# a_6638_19998# VGND.t94 sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.145 ps=1.58 w=0.5 l=20
**devattr s=5800,316 d=5800,316
X171 VAPWR.t19 a_21737_7899.t11 ua[0].t0 VAPWR.t18 sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=8.5 l=1
**devattr s=49300,1758 d=98600,3516
X172 a_7586_26859# a_9886_27155# VGND.t6 sky130_fd_pr__res_xhigh_po_0p35 l=9.5
X173 Timming_0.Vd.t3 a_16597_7688.t42 a_16597_7688.t43 VGND.t50 sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=10 l=0.5
**devattr s=58000,2058 d=58000,2058
X174 a_10404_14647.t8 a_6404_16954.t10 a_6064_20056# VAPWR.t6 sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.87 ps=6.58 w=3 l=20
**devattr s=34800,1316 d=34800,1316
X175 a_6061_11160.t0 COMP_2_0.vin_n.t3 a_5453_6051.t6 VAPWR.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=2.5 l=2.4
**devattr s=29000,1116 d=29000,1116
X176 a_18714_5807# a_19010_2607# VGND.t88 sky130_fd_pr__res_xhigh_po_0p35 l=14
X177 VGND.t100 VGND.t101 VGND.t6 sky130_fd_pr__res_xhigh_po_0p35 l=9.5
X178 VGND.t78 VGND.t79 BIAS_1_0.XQ12.Emitter sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X179 VGND.t29 COMP_2_0.vb.t10 a_10040_19998# VGND.t28 sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.145 ps=1.58 w=0.5 l=20
**devattr s=5800,316 d=5800,316
X180 Timming_0.Vd.t2 a_16597_7688.t24 a_16597_7688.t25 VGND.t112 sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=10 l=0.5
**devattr s=58000,2058 d=58000,2058
X181 a_8279_30718# VGND.t133 a_5450_30348# VAPWR.t12 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=10
**devattr s=11600,516 d=11600,516
X182 a_19306_5807# a_19010_2607# VGND.t99 sky130_fd_pr__res_xhigh_po_0p35 l=14
R0 a_9039_8199.n4 a_9039_8199.t3 95.9785
R1 a_9039_8199.t1 a_9039_8199.n12 95.9785
R2 a_9039_8199.n2 a_9039_8199.t4 91.4057
R3 a_9039_8199.n1 a_9039_8199.t5 27.9381
R4 a_9039_8199.n8 a_9039_8199.t6 27.4879
R5 a_9039_8199.n10 a_9039_8199.t0 27.3045
R6 a_9039_8199.n5 a_9039_8199.t2 27.3045
R7 a_9039_8199.n2 a_9039_8199.n0 5.45874
R8 a_9039_8199.n3 a_9039_8199.n2 3.2055
R9 a_9039_8199.n7 a_9039_8199.n1 1.86015
R10 a_9039_8199.n9 a_9039_8199.n8 1.69168
R11 a_9039_8199.n5 a_9039_8199.n4 1.47566
R12 a_9039_8199.n12 a_9039_8199.n11 1.27624
R13 a_9039_8199.n10 a_9039_8199.n0 0.96686
R14 a_9039_8199.n6 a_9039_8199.n3 0.789175
R15 a_9039_8199.n8 a_9039_8199.n7 0.4575
R16 a_9039_8199.n9 a_9039_8199.n1 0.4345
R17 a_9039_8199.n4 a_9039_8199.n3 0.25257
R18 a_9039_8199.n12 a_9039_8199.n0 0.25257
R19 a_9039_8199.n11 a_9039_8199.n10 0.189054
R20 a_9039_8199.n6 a_9039_8199.n5 0.189054
R21 a_9039_8199.n11 a_9039_8199.n9 0.0222391
R22 a_9039_8199.n7 a_9039_8199.n6 0.0113696
R23 a_9577_9007.n3 a_9577_9007.t1 231.671
R24 a_9577_9007.t0 a_9577_9007.n3 113.957
R25 a_9577_9007.n1 a_9577_9007.t5 100.364
R26 a_9577_9007.n0 a_9577_9007.t4 100.364
R27 a_9577_9007.n1 a_9577_9007.t3 97.7554
R28 a_9577_9007.n0 a_9577_9007.t2 97.7554
R29 a_9577_9007.n3 a_9577_9007.n2 1.91964
R30 a_9577_9007.n2 a_9577_9007.n1 0.995692
R31 a_9577_9007.n2 a_9577_9007.n0 0.995692
R32 VAPWR.n330 VAPWR.n197 6556.97
R33 VAPWR.n277 VAPWR.n236 6556.97
R34 VAPWR.n328 VAPWR.n198 6556.97
R35 VAPWR.n321 VAPWR.n239 6556.97
R36 VAPWR.n290 VAPWR.n261 5413.04
R37 VAPWR.n261 VAPWR.n257 5413.04
R38 VAPWR.n260 VAPWR.n257 5413.04
R39 VAPWR.n290 VAPWR.n260 5413.04
R40 VAPWR.n259 VAPWR.n255 5181.1
R41 VAPWR.n291 VAPWR.n255 5181.1
R42 VAPWR.n291 VAPWR.n254 5181.1
R43 VAPWR.n259 VAPWR.n254 5181.1
R44 VAPWR.n145 VAPWR.n19 4984.55
R45 VAPWR.n145 VAPWR.n20 4984.55
R46 VAPWR.n88 VAPWR.n20 4984.55
R47 VAPWR.n88 VAPWR.n19 4984.55
R48 VAPWR.n212 VAPWR.n211 4689.72
R49 VAPWR.n220 VAPWR.n203 4689.72
R50 VAPWR.n430 VAPWR.n400 4302.52
R51 VAPWR.n430 VAPWR.n401 4302.52
R52 VAPWR.n428 VAPWR.n401 4302.52
R53 VAPWR.n428 VAPWR.n400 4302.52
R54 VAPWR.n235 VAPWR.n198 4251.41
R55 VAPWR.n236 VAPWR.n235 4251.41
R56 VAPWR.n324 VAPWR.n196 4251.41
R57 VAPWR.n324 VAPWR.n323 4251.41
R58 VAPWR.n323 VAPWR.n322 4251.41
R59 VAPWR.n322 VAPWR.n232 4251.41
R60 VAPWR.n238 VAPWR.n197 4251.41
R61 VAPWR.n321 VAPWR.n238 4251.41
R62 VAPWR.n205 VAPWR.n202 4194.41
R63 VAPWR.n206 VAPWR.n205 4194.41
R64 VAPWR.n154 VAPWR.n5 2832.31
R65 VAPWR.n153 VAPWR.n5 2832.31
R66 VAPWR.n154 VAPWR.n6 2832.31
R67 VAPWR.n153 VAPWR.n6 2832.31
R68 VAPWR.n366 VAPWR.n365 2822.48
R69 VAPWR.n350 VAPWR.n349 2822.48
R70 VAPWR.n304 VAPWR.n298 2812.66
R71 VAPWR.n301 VAPWR.n300 2812.66
R72 VAPWR.n173 VAPWR.n171 2310.18
R73 VAPWR.n175 VAPWR.n171 2310.18
R74 VAPWR.n175 VAPWR.n170 2310.18
R75 VAPWR.n173 VAPWR.n170 2310.18
R76 VAPWR.n330 VAPWR.n196 2305.55
R77 VAPWR.n277 VAPWR.n232 2305.55
R78 VAPWR.n328 VAPWR.n196 2305.55
R79 VAPWR.n235 VAPWR.n230 2305.55
R80 VAPWR.n323 VAPWR.n230 2305.55
R81 VAPWR.n323 VAPWR.n231 2305.55
R82 VAPWR.n238 VAPWR.n231 2305.55
R83 VAPWR.n239 VAPWR.n232 2305.55
R84 VAPWR.n358 VAPWR.n347 2285.9
R85 VAPWR.n366 VAPWR.n347 2285.9
R86 VAPWR.n349 VAPWR.n348 2285.9
R87 VAPWR.n361 VAPWR.n348 2285.9
R88 VAPWR.n208 VAPWR.n207 1831.13
R89 VAPWR.n424 VAPWR.n405 1643.17
R90 VAPWR.n404 VAPWR.n403 1643.17
R91 VAPWR.n107 VAPWR.n58 1623.52
R92 VAPWR.n107 VAPWR.n61 1623.52
R93 VAPWR.n80 VAPWR.n61 1623.52
R94 VAPWR.n80 VAPWR.n58 1623.52
R95 VAPWR.n131 VAPWR.n22 1623.52
R96 VAPWR.n131 VAPWR.n23 1623.52
R97 VAPWR.n143 VAPWR.n22 1623.52
R98 VAPWR.n143 VAPWR.n23 1623.52
R99 VAPWR.n125 VAPWR.n44 1623.52
R100 VAPWR.n44 VAPWR.n43 1623.52
R101 VAPWR.n125 VAPWR.n34 1623.52
R102 VAPWR.n43 VAPWR.n34 1623.52
R103 VAPWR.n30 VAPWR.n21 1623.52
R104 VAPWR.n134 VAPWR.n21 1623.52
R105 VAPWR.n134 VAPWR.n133 1623.52
R106 VAPWR.n133 VAPWR.n30 1623.52
R107 VAPWR.n126 VAPWR.n39 1623.52
R108 VAPWR.n42 VAPWR.n39 1623.52
R109 VAPWR.n42 VAPWR.n38 1623.52
R110 VAPWR.n126 VAPWR.n38 1623.52
R111 VAPWR.n109 VAPWR.n60 1623.52
R112 VAPWR.n110 VAPWR.n109 1623.52
R113 VAPWR.n110 VAPWR.n59 1623.52
R114 VAPWR.n60 VAPWR.n59 1623.52
R115 VAPWR.n92 VAPWR.n74 1623.52
R116 VAPWR.n94 VAPWR.n73 1623.52
R117 VAPWR.n94 VAPWR.n74 1623.52
R118 VAPWR.n78 VAPWR.n77 1623.52
R119 VAPWR.n79 VAPWR.n72 1623.52
R120 VAPWR.n79 VAPWR.n78 1623.52
R121 VAPWR.n367 VAPWR.t26 1391.5
R122 VAPWR.n367 VAPWR.t12 1391.5
R123 VAPWR.n359 VAPWR.n350 942.51
R124 VAPWR.n365 VAPWR.n360 942.51
R125 VAPWR.n304 VAPWR.n303 938.761
R126 VAPWR.n302 VAPWR.n301 938.761
R127 VAPWR.n325 VAPWR.n229 814.307
R128 VAPWR.n233 VAPWR.n229 814.307
R129 VAPWR.n216 VAPWR.n201 804.519
R130 VAPWR.n326 VAPWR.n325 803.389
R131 VAPWR.n279 VAPWR.n233 801.13
R132 VAPWR.n222 VAPWR.n201 800.378
R133 VAPWR.t6 VAPWR.n256 792.155
R134 VAPWR.t6 VAPWR.n258 792.155
R135 VAPWR.n287 VAPWR.n286 740.268
R136 VAPWR.n240 VAPWR.n195 722.362
R137 VAPWR.n251 VAPWR.n250 691.201
R138 VAPWR.n286 VAPWR.n253 615.467
R139 VAPWR.n403 VAPWR.n402 556.174
R140 VAPWR.n425 VAPWR.n424 556.174
R141 VAPWR.n368 VAPWR.n347 536.587
R142 VAPWR.n368 VAPWR.n348 536.587
R143 VAPWR.n212 VAPWR.n202 495.31
R144 VAPWR.n220 VAPWR.n202 495.31
R145 VAPWR.n214 VAPWR.n206 495.31
R146 VAPWR.n218 VAPWR.n206 495.31
R147 VAPWR.n266 VAPWR.n229 446.118
R148 VAPWR.n241 VAPWR.n229 446.118
R149 VAPWR.n242 VAPWR.n241 438.589
R150 VAPWR.n267 VAPWR.n266 431.06
R151 VAPWR.n329 VAPWR.t3 411.135
R152 VAPWR.n234 VAPWR.t3 411.135
R153 VAPWR.t1 VAPWR.n234 411.135
R154 VAPWR.t1 VAPWR.n237 411.135
R155 VAPWR.t2 VAPWR.n171 293.449
R156 VAPWR.t31 VAPWR.n170 290.765
R157 VAPWR.n17 VAPWR.n14 254.031
R158 VAPWR.n276 VAPWR.n275 230.196
R159 VAPWR.n159 VAPWR.t25 229.987
R160 VAPWR.n313 VAPWR.t5 229.881
R161 VAPWR.n289 VAPWR.n288 216.928
R162 VAPWR.n208 VAPWR.n200 213.859
R163 VAPWR.t36 VAPWR.t31 212.006
R164 VAPWR.t7 VAPWR.t2 212.006
R165 VAPWR.n180 VAPWR.n179 204.71
R166 VAPWR.n292 VAPWR.n253 203.873
R167 VAPWR.n209 VAPWR.n207 189.806
R168 VAPWR.n269 VAPWR.n268 172.35
R169 VAPWR.n289 VAPWR.n262 166.397
R170 VAPWR.n268 VAPWR.n267 161.91
R171 VAPWR.n267 VAPWR.n265 161.91
R172 VAPWR.n129 VAPWR.n24 140.048
R173 VAPWR.n128 VAPWR.n36 140.048
R174 VAPWR.t13 VAPWR.n7 136.625
R175 VAPWR.n141 VAPWR.n24 136.282
R176 VAPWR.n129 VAPWR.n35 136.282
R177 VAPWR.n36 VAPWR.n25 136.282
R178 VAPWR.n128 VAPWR.n127 136.282
R179 VAPWR.n55 VAPWR.n35 134.4
R180 VAPWR.n127 VAPWR.n37 134.4
R181 VAPWR.t15 VAPWR.n41 122.63
R182 VAPWR.t15 VAPWR.n31 122.63
R183 VAPWR.n132 VAPWR.t0 122.63
R184 VAPWR.n144 VAPWR.t0 122.63
R185 VAPWR.n285 VAPWR.n283 118.442
R186 VAPWR.n147 VAPWR.n17 118.338
R187 VAPWR.t16 VAPWR.n401 115.294
R188 VAPWR.n283 VAPWR.n282 114.121
R189 VAPWR.t18 VAPWR.n426 108.915
R190 VAPWR.n174 VAPWR.t36 107.346
R191 VAPWR.t9 VAPWR.t18 106.844
R192 VAPWR.t38 VAPWR.t9 106.844
R193 VAPWR.t32 VAPWR.t38 106.844
R194 VAPWR.t22 VAPWR.t20 106.844
R195 VAPWR.t20 VAPWR.t34 106.844
R196 VAPWR.t34 VAPWR.t16 106.844
R197 VAPWR.n370 VAPWR.n369 105.412
R198 VAPWR.n174 VAPWR.t7 104.662
R199 VAPWR.n279 VAPWR.n278 102.572
R200 VAPWR.n369 VAPWR.n346 102.025
R201 VAPWR.n363 VAPWR.n345 99.4821
R202 VAPWR.n357 VAPWR.n356 98.6135
R203 VAPWR.t27 VAPWR.n82 97.9161
R204 VAPWR.n81 VAPWR.t28 97.9161
R205 VAPWR.n364 VAPWR.n362 97.0916
R206 VAPWR.n355 VAPWR.n354 96.1993
R207 VAPWR.n427 VAPWR.n398 93.7086
R208 VAPWR.n445 VAPWR.n384 78.8342
R209 VAPWR.n280 VAPWR.n279 77.3125
R210 VAPWR.n318 VAPWR.n246 76.9712
R211 VAPWR.n370 VAPWR.n345 72.6171
R212 VAPWR.n357 VAPWR.n343 71.6805
R213 VAPWR.n362 VAPWR.n346 70.2194
R214 VAPWR.n354 VAPWR.n353 69.3741
R215 VAPWR.n432 VAPWR.n431 67.9353
R216 VAPWR.n145 VAPWR.n144 63.6557
R217 VAPWR.n155 VAPWR.n4 62.248
R218 VAPWR.n441 VAPWR.t30 61.9046
R219 VAPWR.n287 VAPWR.n263 61.3522
R220 VAPWR.n169 VAPWR.n164 59.5526
R221 VAPWR.n172 VAPWR.n167 59.2723
R222 VAPWR.n242 VAPWR.n240 57.5606
R223 VAPWR.n320 VAPWR.n319 56.6292
R224 VAPWR.n135 VAPWR.n29 55.2526
R225 VAPWR.n152 VAPWR.n9 55.06
R226 VAPWR.n213 VAPWR.n211 54.955
R227 VAPWR.n219 VAPWR.n203 54.955
R228 VAPWR.n176 VAPWR.n168 54.8382
R229 VAPWR.n429 VAPWR.t32 53.4225
R230 VAPWR.n429 VAPWR.t22 53.4225
R231 VAPWR.t11 VAPWR.n204 53.012
R232 VAPWR.t14 VAPWR.n204 53.012
R233 VAPWR.n177 VAPWR.n176 52.1671
R234 VAPWR.t24 VAPWR.t28 51.7524
R235 VAPWR.n285 VAPWR.n284 49.9867
R236 VAPWR.n299 VAPWR.n251 48.7693
R237 VAPWR.n157 VAPWR.n3 48.0785
R238 VAPWR.n411 VAPWR.n406 44.0139
R239 VAPWR.n70 VAPWR.n66 43.2599
R240 VAPWR.n319 VAPWR.n318 43.0085
R241 VAPWR.n40 VAPWR.n6 39.8695
R242 VAPWR.n152 VAPWR.n151 39.8173
R243 VAPWR.n132 VAPWR.n31 39.5585
R244 VAPWR.n426 VAPWR.t29 39.3423
R245 VAPWR.n299 VAPWR.n245 39.0126
R246 VAPWR.n41 VAPWR.n40 38.8336
R247 VAPWR.n320 VAPWR.n244 38.2941
R248 VAPWR.n424 VAPWR.n423 37.0005
R249 VAPWR.n403 VAPWR.n385 37.0005
R250 VAPWR.n218 VAPWR.n217 37.0005
R251 VAPWR.n215 VAPWR.n214 37.0005
R252 VAPWR.n221 VAPWR.n220 37.0005
R253 VAPWR.n220 VAPWR.t14 37.0005
R254 VAPWR.n212 VAPWR.n200 37.0005
R255 VAPWR.t11 VAPWR.n212 37.0005
R256 VAPWR.n71 VAPWR.n70 36.2942
R257 VAPWR.n214 VAPWR.n213 36.2812
R258 VAPWR.n219 VAPWR.n218 36.2812
R259 VAPWR.n136 VAPWR.n135 35.2716
R260 VAPWR.n422 VAPWR.n399 35.2005
R261 VAPWR.n104 VAPWR.n103 35.1091
R262 VAPWR.n96 VAPWR.n71 34.5929
R263 VAPWR.n91 VAPWR.n69 34.4978
R264 VAPWR.n136 VAPWR.n28 34.3235
R265 VAPWR.n301 VAPWR.n245 33.9241
R266 VAPWR.n105 VAPWR.n28 33.8494
R267 VAPWR.n70 VAPWR.n63 33.2805
R268 VAPWR.n103 VAPWR.n63 33.2805
R269 VAPWR.n96 VAPWR.n69 32.8916
R270 VAPWR.n105 VAPWR.n104 32.4716
R271 VAPWR.n146 VAPWR.n18 32.0626
R272 VAPWR.t24 VAPWR.n7 31.8521
R273 VAPWR.n40 VAPWR.t13 31.7391
R274 VAPWR.n103 VAPWR.n64 31.3048
R275 VAPWR.n82 VAPWR.n81 30.6143
R276 VAPWR.n410 VAPWR.n407 30.4557
R277 VAPWR.n64 VAPWR.n57 29.7048
R278 VAPWR.n137 VAPWR.n27 29.3391
R279 VAPWR.n395 VAPWR.t17 29.0249
R280 VAPWR.n84 VAPWR.n83 28.8701
R281 VAPWR.n76 VAPWR.n5 28.8395
R282 VAPWR.n388 VAPWR.t19 28.6551
R283 VAPWR.n130 VAPWR.n129 28.6421
R284 VAPWR.n128 VAPWR.n27 28.6421
R285 VAPWR.n83 VAPWR.n57 28.244
R286 VAPWR.n275 VAPWR.n265 27.9958
R287 VAPWR.n422 VAPWR.n421 27.7509
R288 VAPWR.n179 VAPWR.t37 27.6955
R289 VAPWR.n179 VAPWR.t8 27.6955
R290 VAPWR.n130 VAPWR.n33 27.4381
R291 VAPWR.n355 VAPWR.n350 26.4667
R292 VAPWR.n365 VAPWR.n364 26.4505
R293 VAPWR.n305 VAPWR.n304 26.4291
R294 VAPWR.n170 VAPWR.n169 26.4291
R295 VAPWR.n171 VAPWR.n167 26.4291
R296 VAPWR.n15 VAPWR.n6 26.4291
R297 VAPWR.n8 VAPWR.n5 26.4291
R298 VAPWR.n369 VAPWR.n368 26.4291
R299 VAPWR.n368 VAPWR.n367 26.4291
R300 VAPWR.n392 VAPWR.n391 25.7666
R301 VAPWR.n393 VAPWR.n390 25.7666
R302 VAPWR.n394 VAPWR.n389 25.7666
R303 VAPWR.n280 VAPWR.n246 25.2592
R304 VAPWR.n142 VAPWR.n18 24.9717
R305 VAPWR.n84 VAPWR.n45 24.6677
R306 VAPWR.n33 VAPWR.n32 24.5122
R307 VAPWR.n111 VAPWR.n57 24.1783
R308 VAPWR.n293 VAPWR.n250 24.1206
R309 VAPWR.n124 VAPWR.n33 23.994
R310 VAPWR.n97 VAPWR.n68 23.7712
R311 VAPWR.n95 VAPWR.n57 23.1624
R312 VAPWR.n281 VAPWR.n280 23.1556
R313 VAPWR.n90 VAPWR.n84 22.6985
R314 VAPWR.n293 VAPWR.n292 22.5368
R315 VAPWR.n96 VAPWR.n95 22.5021
R316 VAPWR.n222 VAPWR.n221 22.4005
R317 VAPWR.n223 VAPWR.n200 22.2227
R318 VAPWR.n331 VAPWR.n195 22.0785
R319 VAPWR.n142 VAPWR.n141 20.3009
R320 VAPWR.n29 VAPWR.n25 20.3009
R321 VAPWR.n327 VAPWR.n326 19.6
R322 VAPWR.n243 VAPWR.n242 19.0541
R323 VAPWR.n32 VAPWR.n18 18.76
R324 VAPWR.n123 VAPWR.n45 18.6045
R325 VAPWR.n88 VAPWR.n76 18.5122
R326 VAPWR.n124 VAPWR.n123 18.5009
R327 VAPWR.n127 VAPWR.n126 18.5005
R328 VAPWR.n126 VAPWR.t15 18.5005
R329 VAPWR.n42 VAPWR.n28 18.5005
R330 VAPWR.t15 VAPWR.n42 18.5005
R331 VAPWR.n36 VAPWR.n30 18.5005
R332 VAPWR.n30 VAPWR.t0 18.5005
R333 VAPWR.n43 VAPWR.n35 18.5005
R334 VAPWR.t15 VAPWR.n43 18.5005
R335 VAPWR.n24 VAPWR.n23 18.5005
R336 VAPWR.n23 VAPWR.t0 18.5005
R337 VAPWR.n78 VAPWR.n63 18.5005
R338 VAPWR.t27 VAPWR.n78 18.5005
R339 VAPWR.n60 VAPWR.n45 18.5005
R340 VAPWR.n60 VAPWR.t28 18.5005
R341 VAPWR.n92 VAPWR.n91 18.5005
R342 VAPWR.n89 VAPWR.n88 18.5005
R343 VAPWR.n95 VAPWR.n72 18.5005
R344 VAPWR.n111 VAPWR.n58 18.5005
R345 VAPWR.n58 VAPWR.t28 18.5005
R346 VAPWR.n95 VAPWR.n94 18.5005
R347 VAPWR.n94 VAPWR.t27 18.5005
R348 VAPWR.n111 VAPWR.n110 18.5005
R349 VAPWR.n110 VAPWR.t28 18.5005
R350 VAPWR.n104 VAPWR.n61 18.5005
R351 VAPWR.n61 VAPWR.t28 18.5005
R352 VAPWR.n125 VAPWR.n124 18.5005
R353 VAPWR.t15 VAPWR.n125 18.5005
R354 VAPWR.n32 VAPWR.n22 18.5005
R355 VAPWR.n22 VAPWR.t0 18.5005
R356 VAPWR.n135 VAPWR.n134 18.5005
R357 VAPWR.n134 VAPWR.t0 18.5005
R358 VAPWR.n146 VAPWR.n145 18.5005
R359 VAPWR.n112 VAPWR.n111 18.2354
R360 VAPWR.n93 VAPWR.n92 18.1071
R361 VAPWR.n75 VAPWR.n72 18.1071
R362 VAPWR.n418 VAPWR.n417 17.8322
R363 VAPWR.n83 VAPWR.n74 16.8187
R364 VAPWR.n82 VAPWR.n74 16.8187
R365 VAPWR.n83 VAPWR.n59 16.8187
R366 VAPWR.n81 VAPWR.n59 16.8187
R367 VAPWR.n73 VAPWR.n69 16.8187
R368 VAPWR.n77 VAPWR.n71 16.8187
R369 VAPWR.n79 VAPWR.n64 16.8187
R370 VAPWR.n82 VAPWR.n79 16.8187
R371 VAPWR.n80 VAPWR.n64 16.8187
R372 VAPWR.n81 VAPWR.n80 16.8187
R373 VAPWR.n107 VAPWR.n106 16.8187
R374 VAPWR.n108 VAPWR.n107 16.8187
R375 VAPWR.n62 VAPWR.n38 16.8187
R376 VAPWR.n41 VAPWR.n38 16.8187
R377 VAPWR.n54 VAPWR.n44 16.8187
R378 VAPWR.n44 VAPWR.n41 16.8187
R379 VAPWR.n109 VAPWR.n47 16.8187
R380 VAPWR.n109 VAPWR.n108 16.8187
R381 VAPWR.n39 VAPWR.n27 16.8187
R382 VAPWR.n39 VAPWR.n31 16.8187
R383 VAPWR.n133 VAPWR.n27 16.8187
R384 VAPWR.n133 VAPWR.n132 16.8187
R385 VAPWR.n130 VAPWR.n34 16.8187
R386 VAPWR.n34 VAPWR.n31 16.8187
R387 VAPWR.n131 VAPWR.n130 16.8187
R388 VAPWR.n132 VAPWR.n131 16.8187
R389 VAPWR.n29 VAPWR.n21 16.8187
R390 VAPWR.n144 VAPWR.n21 16.8187
R391 VAPWR.n143 VAPWR.n142 16.8187
R392 VAPWR.n144 VAPWR.n143 16.8187
R393 VAPWR.n332 VAPWR.n331 16.5345
R394 VAPWR.n77 VAPWR.n75 16.4611
R395 VAPWR.n93 VAPWR.n73 16.4611
R396 VAPWR.n306 VAPWR.n250 15.5663
R397 VAPWR.n284 VAPWR.n255 15.4172
R398 VAPWR.n258 VAPWR.n255 15.4172
R399 VAPWR.n281 VAPWR.n254 15.4172
R400 VAPWR.n256 VAPWR.n254 15.4172
R401 VAPWR.n173 VAPWR.n172 15.4172
R402 VAPWR.n174 VAPWR.n173 15.4172
R403 VAPWR.n176 VAPWR.n175 15.4172
R404 VAPWR.n175 VAPWR.n174 15.4172
R405 VAPWR.n228 VAPWR.n227 14.5783
R406 VAPWR.n280 VAPWR.n245 14.4721
R407 VAPWR.n420 VAPWR.n419 14.3877
R408 VAPWR.n327 VAPWR.n228 14.105
R409 VAPWR.n16 VAPWR.n15 13.4801
R410 VAPWR.n423 VAPWR.n422 12.4179
R411 VAPWR.n410 VAPWR.n404 12.3338
R412 VAPWR.n421 VAPWR.n405 12.3338
R413 VAPWR.n269 VAPWR.n228 12.1251
R414 VAPWR.n288 VAPWR.n261 11.7128
R415 VAPWR.n261 VAPWR.n258 11.563
R416 VAPWR.n262 VAPWR.n260 11.563
R417 VAPWR.n260 VAPWR.n256 11.563
R418 VAPWR.n87 VAPWR.n9 11.4968
R419 VAPWR.n90 VAPWR.n89 11.3783
R420 VAPWR.n376 VAPWR 10.6062
R421 VAPWR.n282 VAPWR.n281 10.4866
R422 VAPWR.n16 VAPWR.n10 10.0646
R423 VAPWR.n411 VAPWR.n410 9.71084
R424 VAPWR.n276 VAPWR.n262 9.38472
R425 VAPWR.n420 VAPWR.n387 9.3005
R426 VAPWR.n415 VAPWR.n407 9.3005
R427 VAPWR.n412 VAPWR.n411 9.3005
R428 VAPWR.n224 VAPWR.n223 9.3005
R429 VAPWR.n184 VAPWR.n164 9.3005
R430 VAPWR.n122 VAPWR.n121 9.3005
R431 VAPWR.n372 VAPWR.n371 9.3005
R432 VAPWR.n151 VAPWR.n10 9.28294
R433 VAPWR.n319 VAPWR.n245 9.02171
R434 VAPWR.n9 VAPWR.n8 8.74717
R435 VAPWR.n129 VAPWR.n128 8.74505
R436 VAPWR.n421 VAPWR.n420 8.6533
R437 VAPWR.n431 VAPWR.n399 8.34833
R438 VAPWR.n425 VAPWR.n404 8.09902
R439 VAPWR.n405 VAPWR.n402 8.09902
R440 VAPWR.n274 VAPWR.n270 7.38601
R441 VAPWR.n445 VAPWR.n444 7.06871
R442 VAPWR.n156 VAPWR.n155 6.48
R443 VAPWR.n419 VAPWR.n400 6.37981
R444 VAPWR.n426 VAPWR.n400 6.37981
R445 VAPWR.n401 VAPWR.n398 6.37981
R446 VAPWR.n318 VAPWR.n317 6.27883
R447 VAPWR.n215 VAPWR.n207 6.20324
R448 VAPWR.n419 VAPWR.n418 6.1445
R449 VAPWR.n278 VAPWR.n276 6.05917
R450 VAPWR.n210 VAPWR.n208 6.03479
R451 VAPWR.n17 VAPWR.n16 5.8631
R452 VAPWR.n431 VAPWR.n430 5.78175
R453 VAPWR.n430 VAPWR.n429 5.78175
R454 VAPWR.n428 VAPWR.n427 5.78175
R455 VAPWR.n429 VAPWR.n428 5.78175
R456 VAPWR.n298 VAPWR.n297 5.78175
R457 VAPWR.n300 VAPWR.n299 5.78175
R458 VAPWR.n153 VAPWR.n152 5.78175
R459 VAPWR.t24 VAPWR.n153 5.78175
R460 VAPWR.n155 VAPWR.n154 5.78175
R461 VAPWR.n154 VAPWR.t24 5.78175
R462 VAPWR.n358 VAPWR.n357 5.78175
R463 VAPWR.n366 VAPWR.n345 5.78175
R464 VAPWR.t12 VAPWR.n366 5.78175
R465 VAPWR.n362 VAPWR.n361 5.78175
R466 VAPWR.n354 VAPWR.n349 5.78175
R467 VAPWR.t26 VAPWR.n349 5.78175
R468 VAPWR.n328 VAPWR.n327 5.60656
R469 VAPWR.n329 VAPWR.n328 5.60656
R470 VAPWR.n331 VAPWR.n330 5.60656
R471 VAPWR.n330 VAPWR.n329 5.60656
R472 VAPWR.n266 VAPWR.n230 5.60656
R473 VAPWR.n234 VAPWR.n230 5.60656
R474 VAPWR.n241 VAPWR.n231 5.60656
R475 VAPWR.n234 VAPWR.n231 5.60656
R476 VAPWR.n278 VAPWR.n277 5.60656
R477 VAPWR.n277 VAPWR.n237 5.60656
R478 VAPWR.n246 VAPWR.n239 5.60656
R479 VAPWR.n239 VAPWR.n237 5.60656
R480 VAPWR.n210 VAPWR.n209 5.57764
R481 VAPWR.n216 VAPWR.n215 5.52379
R482 VAPWR.n217 VAPWR.n216 5.52379
R483 VAPWR.n273 VAPWR.n272 5.33984
R484 VAPWR.n414 VAPWR.n413 4.90422
R485 VAPWR.n122 VAPWR.n47 4.86113
R486 VAPWR.n423 VAPWR.n406 4.8005
R487 VAPWR.n108 VAPWR.n7 4.77187
R488 VAPWR.n55 VAPWR.n54 4.76623
R489 VAPWR.n62 VAPWR.n37 4.76623
R490 VAPWR.n280 VAPWR.n252 4.71845
R491 VAPWR.n106 VAPWR.n105 4.65025
R492 VAPWR.n217 VAPWR.n195 4.64707
R493 VAPWR.n177 VAPWR.n167 4.62502
R494 VAPWR.n297 VAPWR.n296 4.59537
R495 VAPWR.n140 VAPWR.n25 4.58155
R496 VAPWR.n336 VAPWR.n335 4.501
R497 VAPWR.n439 VAPWR.n387 4.5005
R498 VAPWR.n310 VAPWR.n309 4.5005
R499 VAPWR.n311 VAPWR.n248 4.5005
R500 VAPWR.n182 VAPWR.n181 4.5005
R501 VAPWR.n185 VAPWR.n184 4.5005
R502 VAPWR.n99 VAPWR.n66 4.5005
R503 VAPWR.n101 VAPWR.n100 4.5005
R504 VAPWR.t29 VAPWR.n402 4.17553
R505 VAPWR.t29 VAPWR.n425 4.17553
R506 VAPWR.n169 VAPWR.n168 4.04695
R507 VAPWR.n292 VAPWR.n291 3.99394
R508 VAPWR.n302 VAPWR.n298 3.84478
R509 VAPWR.n303 VAPWR.n300 3.84478
R510 VAPWR.n359 VAPWR.n358 3.84385
R511 VAPWR.n361 VAPWR.n360 3.84385
R512 VAPWR.n46 VAPWR.n20 3.70808
R513 VAPWR.n221 VAPWR.n199 3.46717
R514 VAPWR.n338 VAPWR.n188 3.43119
R515 VAPWR.n337 VAPWR.n189 3.4105
R516 VAPWR.n189 VAPWR.n188 3.4105
R517 VAPWR.n391 VAPWR.t10 3.25874
R518 VAPWR.n391 VAPWR.t39 3.25874
R519 VAPWR.n390 VAPWR.t33 3.25874
R520 VAPWR.n390 VAPWR.t23 3.25874
R521 VAPWR.n389 VAPWR.t21 3.25874
R522 VAPWR.n389 VAPWR.t35 3.25874
R523 VAPWR.t27 VAPWR.n76 3.13387
R524 VAPWR.n286 VAPWR.n285 3.13299
R525 VAPWR.n290 VAPWR.n289 3.03329
R526 VAPWR.t6 VAPWR.n290 3.03329
R527 VAPWR.n283 VAPWR.n259 3.03329
R528 VAPWR.t6 VAPWR.n259 3.03329
R529 VAPWR.n283 VAPWR.n257 3.03329
R530 VAPWR.t6 VAPWR.n257 3.03329
R531 VAPWR.n291 VAPWR.t6 3.03329
R532 VAPWR.n321 VAPWR.n320 3.03329
R533 VAPWR.t1 VAPWR.n321 3.03329
R534 VAPWR.n240 VAPWR.n197 3.03329
R535 VAPWR.t3 VAPWR.n197 3.03329
R536 VAPWR.n211 VAPWR.n210 3.03329
R537 VAPWR.n205 VAPWR.n201 3.03329
R538 VAPWR.n205 VAPWR.n204 3.03329
R539 VAPWR.n203 VAPWR.n194 3.03329
R540 VAPWR.n265 VAPWR.n236 3.03329
R541 VAPWR.t1 VAPWR.n236 3.03329
R542 VAPWR.n268 VAPWR.n198 3.03329
R543 VAPWR.n198 VAPWR.t3 3.03329
R544 VAPWR.n322 VAPWR.n233 3.03329
R545 VAPWR.n322 VAPWR.t1 3.03329
R546 VAPWR.n325 VAPWR.n324 3.03329
R547 VAPWR.n324 VAPWR.t3 3.03329
R548 VAPWR.n19 VAPWR.n10 3.03329
R549 VAPWR.t13 VAPWR.n19 3.03329
R550 VAPWR.t13 VAPWR.n20 3.03329
R551 VAPWR.n448 VAPWR.n381 2.76526
R552 VAPWR.n272 VAPWR.n249 2.73361
R553 VAPWR.n282 VAPWR.n264 2.53479
R554 VAPWR.n224 VAPWR.n191 2.35179
R555 VAPWR.n285 VAPWR.n263 2.09705
R556 VAPWR.n326 VAPWR.n194 2.07133
R557 VAPWR.n91 VAPWR.n90 2.03902
R558 VAPWR.n417 VAPWR.n407 2.03084
R559 VAPWR.n317 VAPWR.n245 1.9716
R560 VAPWR.n297 VAPWR.n252 1.96973
R561 VAPWR.t12 VAPWR.n360 1.93153
R562 VAPWR.t26 VAPWR.n359 1.93153
R563 VAPWR.t4 VAPWR.n302 1.93057
R564 VAPWR.n303 VAPWR.t4 1.93057
R565 VAPWR.n335 VAPWR.n191 1.89315
R566 VAPWR.n118 VAPWR.n26 1.85564
R567 VAPWR.n372 VAPWR.n344 1.78482
R568 VAPWR.n351 VAPWR.n344 1.78482
R569 VAPWR.n342 VAPWR.n341 1.76185
R570 VAPWR.n117 VAPWR.n116 1.7485
R571 VAPWR.n336 VAPWR.n190 1.74586
R572 VAPWR.n312 VAPWR.n311 1.73031
R573 VAPWR.n288 VAPWR.n287 1.72305
R574 VAPWR.n432 VAPWR.n398 1.72202
R575 VAPWR.n116 VAPWR.n51 1.69007
R576 VAPWR.n274 VAPWR.n273 1.67948
R577 VAPWR.n50 VAPWR.n26 1.65581
R578 VAPWR.n141 VAPWR.n140 1.61734
R579 VAPWR.n376 VAPWR 1.58252
R580 VAPWR.n114 VAPWR.n53 1.56843
R581 VAPWR.n187 VAPWR.n160 1.45744
R582 VAPWR.n139 VAPWR.n138 1.44157
R583 VAPWR.n165 VAPWR.n164 1.40196
R584 VAPWR.n334 VAPWR.n192 1.32787
R585 VAPWR.n296 VAPWR.n293 1.28597
R586 VAPWR.n375 VAPWR.n341 1.26013
R587 VAPWR.n98 VAPWR.n67 1.21343
R588 VAPWR.n413 VAPWR.n382 1.19878
R589 VAPWR.n49 VAPWR.n13 1.18185
R590 VAPWR.n270 VAPWR.n269 1.16893
R591 VAPWR.n435 VAPWR.n434 1.14155
R592 VAPWR.n276 VAPWR.n264 1.13909
R593 VAPWR.n15 VAPWR.n14 1.13324
R594 VAPWR.n150 VAPWR.n11 1.09704
R595 VAPWR.n180 VAPWR.n178 0.99906
R596 VAPWR.n439 VAPWR.n438 0.997283
R597 VAPWR.n332 VAPWR.n194 0.99515
R598 VAPWR.n99 VAPWR.n98 0.993269
R599 VAPWR.n433 VAPWR.n380 0.94407
R600 VAPWR.n315 VAPWR.n248 0.943921
R601 VAPWR.n381 VAPWR.n380 0.928345
R602 VAPWR.n97 VAPWR.n65 0.917167
R603 VAPWR.n68 VAPWR.n52 0.902702
R604 VAPWR.n187 VAPWR.n186 0.881527
R605 VAPWR.n442 VAPWR.n382 0.881314
R606 VAPWR.n438 VAPWR.n396 0.874399
R607 VAPWR.n437 VAPWR.n436 0.867309
R608 VAPWR.n364 VAPWR.n363 0.852922
R609 VAPWR.n188 VAPWR.n187 0.848609
R610 VAPWR.n379 VAPWR 0.84274
R611 VAPWR.n118 VAPWR.n117 0.841629
R612 VAPWR.n408 VAPWR.n386 0.836361
R613 VAPWR.n433 VAPWR.n383 0.816018
R614 VAPWR.n123 VAPWR.n122 0.812362
R615 VAPWR.n371 VAPWR.n370 0.812207
R616 VAPWR.n392 VAPWR.n388 0.809067
R617 VAPWR.n100 VAPWR.n99 0.807718
R618 VAPWR.n149 VAPWR.n148 0.805975
R619 VAPWR.n112 VAPWR.n37 0.801818
R620 VAPWR.n227 VAPWR.n199 0.8005
R621 VAPWR.n352 VAPWR.n346 0.785406
R622 VAPWR.n451 VAPWR 0.777997
R623 VAPWR.n409 VAPWR.n406 0.7755
R624 VAPWR.n374 VAPWR.n373 0.77267
R625 VAPWR.n356 VAPWR.n355 0.76856
R626 VAPWR.n101 VAPWR.n65 0.76771
R627 VAPWR.n172 VAPWR.n166 0.747945
R628 VAPWR.n115 VAPWR.n52 0.747335
R629 VAPWR.n182 VAPWR.n178 0.732569
R630 VAPWR.n315 VAPWR.n314 0.728797
R631 VAPWR.n12 VAPWR.n2 0.705003
R632 VAPWR.n409 VAPWR.n397 0.689864
R633 VAPWR.n379 VAPWR.n378 0.683528
R634 VAPWR.n184 VAPWR.n163 0.675345
R635 VAPWR.n120 VAPWR.n119 0.671929
R636 VAPWR.n147 VAPWR.n146 0.670267
R637 VAPWR.n284 VAPWR.n253 0.662569
R638 VAPWR.n356 VAPWR.n342 0.629958
R639 VAPWR.n182 VAPWR.n166 0.6205
R640 VAPWR.n183 VAPWR.n165 0.6205
R641 VAPWR.n363 VAPWR.n344 0.609139
R642 VAPWR.n178 VAPWR.n177 0.58175
R643 VAPWR.n168 VAPWR.n163 0.58175
R644 VAPWR.n443 VAPWR.n386 0.565798
R645 VAPWR.n375 VAPWR.n374 0.558331
R646 VAPWR.n163 VAPWR.n161 0.527844
R647 VAPWR.n412 VAPWR.n409 0.521249
R648 VAPWR.n103 VAPWR.n102 0.518863
R649 VAPWR.n139 VAPWR.n13 0.514931
R650 VAPWR.n8 VAPWR.n3 0.498278
R651 VAPWR.n158 VAPWR.n1 0.492548
R652 VAPWR.n418 VAPWR.n385 0.475674
R653 VAPWR.n427 VAPWR.n384 0.453025
R654 VAPWR.n393 VAPWR.n392 0.439276
R655 VAPWR.n394 VAPWR.n393 0.439276
R656 VAPWR.n395 VAPWR.n394 0.439276
R657 VAPWR.t14 VAPWR.n219 0.434565
R658 VAPWR.n213 VAPWR.t11 0.434565
R659 VAPWR.n148 VAPWR.n147 0.423227
R660 VAPWR.n334 VAPWR.n333 0.41025
R661 VAPWR.n415 VAPWR.n414 0.392464
R662 VAPWR.n12 VAPWR.n4 0.390448
R663 VAPWR.n307 VAPWR.n306 0.388
R664 VAPWR.n444 VAPWR.n385 0.386579
R665 VAPWR.n333 VAPWR.n193 0.382248
R666 VAPWR.n56 VAPWR.n55 0.380072
R667 VAPWR.n52 VAPWR.n48 0.370966
R668 VAPWR.n225 VAPWR.n199 0.358192
R669 VAPWR.n227 VAPWR.n226 0.358192
R670 VAPWR.n440 VAPWR.n388 0.331455
R671 VAPWR.n148 VAPWR.n13 0.330762
R672 VAPWR.n97 VAPWR.n96 0.325103
R673 VAPWR.n138 VAPWR.n137 0.32119
R674 VAPWR.n306 VAPWR.n305 0.300969
R675 VAPWR.n314 VAPWR.n313 0.3005
R676 VAPWR.n443 VAPWR.n387 0.28722
R677 VAPWR.n183 VAPWR.n162 0.28175
R678 VAPWR.n106 VAPWR.n62 0.264091
R679 VAPWR.n313 VAPWR.n312 0.259711
R680 VAPWR.n335 VAPWR.n334 0.255999
R681 VAPWR.n67 VAPWR.n0 0.255814
R682 VAPWR.n225 VAPWR.n224 0.253086
R683 VAPWR.n434 VAPWR.n433 0.245398
R684 VAPWR.n113 VAPWR.n112 0.23246
R685 VAPWR.n156 VAPWR.n2 0.227329
R686 VAPWR.n442 VAPWR.n441 0.222032
R687 VAPWR.n186 VAPWR.n185 0.221874
R688 VAPWR.n374 VAPWR.n342 0.219746
R689 VAPWR.n150 VAPWR.n149 0.216251
R690 VAPWR.n89 VAPWR.n87 0.213833
R691 VAPWR.n244 VAPWR.n243 0.21339
R692 VAPWR.n186 VAPWR.n161 0.206607
R693 VAPWR.n273 VAPWR.n271 0.20095
R694 VAPWR.n450 VAPWR.n449 0.195357
R695 VAPWR.n137 VAPWR.n136 0.190599
R696 VAPWR.n54 VAPWR.n47 0.190286
R697 VAPWR.n271 VAPWR.n247 0.190172
R698 VAPWR.t27 VAPWR.n93 0.188563
R699 VAPWR.t27 VAPWR.n75 0.188563
R700 VAPWR.n223 VAPWR.n222 0.178278
R701 VAPWR.n307 VAPWR.n249 0.176839
R702 VAPWR.n160 VAPWR.n159 0.176252
R703 VAPWR.n444 VAPWR.n443 0.172722
R704 VAPWR.n114 VAPWR.n113 0.172722
R705 VAPWR.n56 VAPWR.n50 0.172722
R706 VAPWR.n149 VAPWR.n12 0.171703
R707 VAPWR.n3 VAPWR.n1 0.166571
R708 VAPWR.n435 VAPWR.n396 0.15931
R709 VAPWR.n161 VAPWR 0.158897
R710 VAPWR.n121 VAPWR.n120 0.15335
R711 VAPWR.n226 VAPWR.n193 0.153086
R712 VAPWR.n123 VAPWR.n46 0.148111
R713 VAPWR.n434 VAPWR.n384 0.141409
R714 VAPWR.n272 VAPWR.n263 0.141409
R715 VAPWR.n353 VAPWR.n341 0.139306
R716 VAPWR.n352 VAPWR.n351 0.139306
R717 VAPWR.n417 VAPWR.n416 0.137265
R718 VAPWR.n121 VAPWR.n48 0.135863
R719 VAPWR VAPWR.n451 0.13369
R720 VAPWR.n312 VAPWR 0.12886
R721 VAPWR.n371 VAPWR.n343 0.125378
R722 VAPWR.n270 VAPWR.n193 0.124924
R723 VAPWR.n87 VAPWR.n86 0.121279
R724 VAPWR.n160 VAPWR.n0 0.121252
R725 VAPWR.n305 VAPWR.n251 0.120688
R726 VAPWR.n140 VAPWR.n139 0.115315
R727 VAPWR.n86 VAPWR.n68 0.115063
R728 VAPWR.n317 VAPWR.n316 0.106182
R729 VAPWR.n396 VAPWR.n395 0.105092
R730 VAPWR.n446 VAPWR.n445 0.095398
R731 VAPWR.n340 VAPWR.n339 0.0952222
R732 VAPWR.n166 VAPWR.n165 0.0939307
R733 VAPWR.n11 VAPWR.n1 0.0929757
R734 VAPWR.n338 VAPWR.n337 0.0928461
R735 VAPWR.n378 VAPWR 0.0919292
R736 VAPWR.n381 VAPWR 0.0897857
R737 VAPWR.n294 VAPWR.n247 0.0857519
R738 VAPWR.n316 VAPWR.n315 0.0841551
R739 VAPWR VAPWR.n375 0.0809707
R740 VAPWR.n386 VAPWR.n383 0.0802354
R741 VAPWR.n157 VAPWR.n156 0.0800031
R742 VAPWR.n209 VAPWR.n191 0.0767295
R743 VAPWR.n158 VAPWR.n157 0.0761098
R744 VAPWR.n443 VAPWR.n442 0.0755
R745 VAPWR.n119 VAPWR.n118 0.0755
R746 VAPWR.n53 VAPWR.n51 0.0755
R747 VAPWR.n98 VAPWR.n97 0.0755
R748 VAPWR.n314 VAPWR.n307 0.0747925
R749 VAPWR.n116 VAPWR.n115 0.0730806
R750 VAPWR.n86 VAPWR.n85 0.0716165
R751 VAPWR.n447 VAPWR.n382 0.0707609
R752 VAPWR.n373 VAPWR.n343 0.069903
R753 VAPWR.n48 VAPWR.n46 0.0678913
R754 VAPWR.n0 VAPWR 0.0664643
R755 VAPWR.n295 VAPWR.n294 0.0655054
R756 VAPWR.n296 VAPWR.n295 0.0650833
R757 VAPWR.n353 VAPWR.n352 0.0608774
R758 VAPWR.n66 VAPWR.n65 0.0607837
R759 VAPWR.n399 VAPWR.n397 0.0601154
R760 VAPWR.n413 VAPWR.n408 0.0597105
R761 VAPWR.n120 VAPWR.n49 0.0574948
R762 VAPWR.n14 VAPWR.n4 0.0556815
R763 VAPWR.n85 VAPWR.n11 0.0492864
R764 VAPWR.n243 VAPWR.n192 0.0491911
R765 VAPWR.n448 VAPWR.n447 0.0491111
R766 VAPWR.n117 VAPWR.n49 0.0481103
R767 VAPWR.n316 VAPWR.n247 0.0460277
R768 VAPWR.n151 VAPWR.n150 0.0454275
R769 VAPWR.n113 VAPWR.n56 0.0426746
R770 VAPWR.n295 VAPWR.n249 0.0403158
R771 VAPWR.n447 VAPWR.n446 0.038
R772 VAPWR.n441 VAPWR.n440 0.0355985
R773 VAPWR.n440 VAPWR.n439 0.0355985
R774 VAPWR.n436 VAPWR.n432 0.0346912
R775 VAPWR.n377 VAPWR.n340 0.0324752
R776 VAPWR.n438 VAPWR.n437 0.0266628
R777 VAPWR.n271 VAPWR.n264 0.0261198
R778 VAPWR.n85 VAPWR.n67 0.0252253
R779 VAPWR.n159 VAPWR.n158 0.0249565
R780 VAPWR.n275 VAPWR.n274 0.0244691
R781 VAPWR.n337 VAPWR.n336 0.0239375
R782 VAPWR.n339 VAPWR.n189 0.0215512
R783 VAPWR.n416 VAPWR.n415 0.0210357
R784 VAPWR.n449 VAPWR.n380 0.0167037
R785 VAPWR.n333 VAPWR.n332 0.0157459
R786 VAPWR.n184 VAPWR.n183 0.0157439
R787 VAPWR.n115 VAPWR.n114 0.0155316
R788 VAPWR.n437 VAPWR.n397 0.0150985
R789 VAPWR.n185 VAPWR.n162 0.014813
R790 VAPWR.n416 VAPWR.n408 0.0147857
R791 VAPWR.n414 VAPWR.n412 0.0147857
R792 VAPWR.n138 VAPWR.n26 0.0145086
R793 VAPWR.n119 VAPWR.n50 0.0140714
R794 VAPWR.n294 VAPWR.n252 0.00892391
R795 VAPWR.n308 VAPWR.n244 0.00861518
R796 VAPWR.n226 VAPWR.n225 0.00825862
R797 VAPWR.n181 VAPWR.n180 0.00810712
R798 VAPWR.n436 VAPWR.n435 0.0062658
R799 VAPWR.n450 VAPWR.n379 0.00605546
R800 VAPWR.n451 VAPWR.n450 0.00603533
R801 VAPWR.n102 VAPWR.n101 0.00457722
R802 VAPWR.n100 VAPWR.n51 0.00402113
R803 VAPWR.n192 VAPWR.n190 0.00349003
R804 VAPWR.n449 VAPWR.n448 0.00296914
R805 VAPWR.n311 VAPWR.n310 0.00257039
R806 VAPWR.n309 VAPWR.n308 0.00234211
R807 VAPWR.n377 VAPWR.n376 0.00220448
R808 VAPWR.n378 VAPWR.n377 0.00219744
R809 VAPWR.n373 VAPWR.n372 0.00176904
R810 VAPWR.n339 VAPWR.n338 0.00156237
R811 VAPWR.n183 VAPWR.n182 0.00151626
R812 VAPWR.n181 VAPWR.n162 0.0014542
R813 VAPWR.n158 VAPWR.n2 0.00128864
R814 VAPWR.n351 VAPWR.n341 0.00113452
R815 VAPWR.n102 VAPWR.n53 0.00104503
R816 VAPWR.n446 VAPWR.n383 0.0010428
R817 VAPWR.n309 VAPWR.n192 0.000763158
R818 VAPWR.n308 VAPWR.n248 0.000763158
R819 VAPWR.n310 VAPWR.n190 0.000758799
R820 VAPWR.n340 VAPWR.n188 0.000594758
R821 VGND.n3269 VGND.n16 561825
R822 VGND.n3144 VGND.n3143 257164
R823 VGND.n3270 VGND.n3269 155264
R824 VGND.n1599 VGND.n1568 39668.3
R825 VGND.n946 VGND.n153 23453.8
R826 VGND.n3104 VGND.n197 18309.4
R827 VGND.n3078 VGND.n222 18309.4
R828 VGND.n1158 VGND.n1089 18309.4
R829 VGND.n3072 VGND.n231 18309.4
R830 VGND.n1090 VGND.n197 17451.9
R831 VGND.n1124 VGND.n1121 17451.9
R832 VGND.n1124 VGND.n198 17451.9
R833 VGND.n1113 VGND.n202 17451.9
R834 VGND.n3099 VGND.n202 17451.9
R835 VGND.n1106 VGND.n1102 17451.9
R836 VGND.n1106 VGND.n203 17451.9
R837 VGND.n1097 VGND.n1096 17451.9
R838 VGND.n1097 VGND.n206 17451.9
R839 VGND.n259 VGND.n210 17451.9
R840 VGND.n3090 VGND.n210 17451.9
R841 VGND.n255 VGND.n251 17451.9
R842 VGND.n255 VGND.n211 17451.9
R843 VGND.n244 VGND.n241 17451.9
R844 VGND.n244 VGND.n214 17451.9
R845 VGND.n235 VGND.n218 17451.9
R846 VGND.n3081 VGND.n218 17451.9
R847 VGND.n3065 VGND.n226 17451.9
R848 VGND.n3065 VGND.n219 17451.9
R849 VGND.n3067 VGND.n230 17451.9
R850 VGND.n3067 VGND.n226 17451.9
R851 VGND.n237 VGND.n233 17451.9
R852 VGND.n237 VGND.n235 17451.9
R853 VGND.n246 VGND.n243 17451.9
R854 VGND.n246 VGND.n241 17451.9
R855 VGND.n253 VGND.n249 17451.9
R856 VGND.n253 VGND.n251 17451.9
R857 VGND.n263 VGND.n261 17451.9
R858 VGND.n263 VGND.n259 17451.9
R859 VGND.n1099 VGND.n1094 17451.9
R860 VGND.n1099 VGND.n1096 17451.9
R861 VGND.n1108 VGND.n1104 17451.9
R862 VGND.n1108 VGND.n1102 17451.9
R863 VGND.n1115 VGND.n1111 17451.9
R864 VGND.n1115 VGND.n1113 17451.9
R865 VGND.n1126 VGND.n1123 17451.9
R866 VGND.n1126 VGND.n1121 17451.9
R867 VGND.n1158 VGND.n1090 17451.9
R868 VGND.n231 VGND.n227 17451.9
R869 VGND.n227 VGND.n222 17451.9
R870 VGND.n1388 VGND.n1313 12805
R871 VGND.n3271 VGND.n15 12805
R872 VGND.n1533 VGND.n1309 12805
R873 VGND.n1496 VGND.n1495 12805
R874 VGND.n3143 VGND.n153 12364
R875 VGND.n1388 VGND.n1387 11947.5
R876 VGND.n1471 VGND.n1316 11947.5
R877 VGND.n1472 VGND.n1471 11947.5
R878 VGND.n1526 VGND.n1320 11947.5
R879 VGND.n1473 VGND.n1320 11947.5
R880 VGND.n1374 VGND.n1322 11947.5
R881 VGND.n1374 VGND.n1373 11947.5
R882 VGND.n1481 VGND.n1342 11947.5
R883 VGND.n1482 VGND.n1481 11947.5
R884 VGND.n1513 VGND.n1346 11947.5
R885 VGND.n1483 VGND.n1346 11947.5
R886 VGND.n1368 VGND.n1348 11947.5
R887 VGND.n1369 VGND.n1368 11947.5
R888 VGND.n3271 VGND.n14 11947.5
R889 VGND.n1507 VGND.n1356 11947.5
R890 VGND.n1507 VGND.n1348 11947.5
R891 VGND.n1355 VGND.n1347 11947.5
R892 VGND.n1513 VGND.n1347 11947.5
R893 VGND.n1518 VGND.n1338 11947.5
R894 VGND.n1518 VGND.n1342 11947.5
R895 VGND.n1335 VGND.n1330 11947.5
R896 VGND.n1335 VGND.n1322 11947.5
R897 VGND.n1329 VGND.n1321 11947.5
R898 VGND.n1526 VGND.n1321 11947.5
R899 VGND.n1531 VGND.n1310 11947.5
R900 VGND.n1531 VGND.n1316 11947.5
R901 VGND.n1387 VGND.n1309 11947.5
R902 VGND.n1502 VGND.n1501 11947.5
R903 VGND.n1501 VGND.n1366 11947.5
R904 VGND.n1489 VGND.n1366 11947.5
R905 VGND.n1489 VGND.n1370 11947.5
R906 VGND.n1496 VGND.n14 11947.5
R907 VGND.n1562 VGND.n1275 11935.9
R908 VGND.n1561 VGND.n1275 11935.9
R909 VGND.n1546 VGND.n1298 11935.9
R910 VGND.n1547 VGND.n1298 11935.9
R911 VGND.n1292 VGND.n1288 11078.4
R912 VGND.n1292 VGND.n1284 11078.4
R913 VGND.n1285 VGND.n1276 11078.4
R914 VGND.n1285 VGND.n1279 11078.4
R915 VGND.n1299 VGND.n1291 11078.4
R916 VGND.n1299 VGND.n1295 11078.4
R917 VGND.n1461 VGND.n1270 9997.86
R918 VGND.n1461 VGND.n1271 9997.86
R919 VGND.n1566 VGND.n1271 9997.86
R920 VGND.n1566 VGND.n1270 9997.86
R921 VGND.n152 VGND.n151 9968.01
R922 VGND.n1568 VGND.n1160 9640.17
R923 VGND.n945 VGND.n298 9328.53
R924 VGND.n943 VGND.n938 9328.53
R925 VGND.n3033 VGND.n278 9328.53
R926 VGND.n802 VGND.n799 9328.53
R927 VGND.n957 VGND.n948 9309.6
R928 VGND.n2598 VGND.n948 9309.6
R929 VGND.n957 VGND.n949 9309.6
R930 VGND.n2598 VGND.n949 9309.6
R931 VGND.n1597 VGND.n1577 9309.6
R932 VGND.n1577 VGND.n716 9309.6
R933 VGND.n1597 VGND.n1578 9309.6
R934 VGND.n1578 VGND.n716 9309.6
R935 VGND.n1569 VGND.n717 8650.98
R936 VGND.n2681 VGND.n717 8650.98
R937 VGND.n1569 VGND.n718 8650.98
R938 VGND.n2681 VGND.n718 8650.98
R939 VGND.n2581 VGND.n955 8650.98
R940 VGND.n2585 VGND.n955 8650.98
R941 VGND.n2585 VGND.n2584 8650.98
R942 VGND.n2584 VGND.n2581 8650.98
R943 VGND.n945 VGND.n944 8569.5
R944 VGND.n944 VGND.n943 8569.5
R945 VGND.n855 VGND.n854 8569.5
R946 VGND.n857 VGND.n855 8569.5
R947 VGND.n936 VGND.n857 8569.5
R948 VGND.n937 VGND.n936 8569.5
R949 VGND.n853 VGND.n852 8569.5
R950 VGND.n863 VGND.n853 8569.5
R951 VGND.n930 VGND.n863 8569.5
R952 VGND.n930 VGND.n929 8569.5
R953 VGND.n851 VGND.n850 8569.5
R954 VGND.n865 VGND.n851 8569.5
R955 VGND.n926 VGND.n865 8569.5
R956 VGND.n927 VGND.n926 8569.5
R957 VGND.n849 VGND.n848 8569.5
R958 VGND.n917 VGND.n849 8569.5
R959 VGND.n918 VGND.n917 8569.5
R960 VGND.n919 VGND.n918 8569.5
R961 VGND.n847 VGND.n846 8569.5
R962 VGND.n872 VGND.n847 8569.5
R963 VGND.n915 VGND.n872 8569.5
R964 VGND.n916 VGND.n915 8569.5
R965 VGND.n845 VGND.n844 8569.5
R966 VGND.n896 VGND.n845 8569.5
R967 VGND.n897 VGND.n896 8569.5
R968 VGND.n898 VGND.n897 8569.5
R969 VGND.n843 VGND.n842 8569.5
R970 VGND.n890 VGND.n843 8569.5
R971 VGND.n891 VGND.n890 8569.5
R972 VGND.n892 VGND.n891 8569.5
R973 VGND.n841 VGND.n840 8569.5
R974 VGND.n889 VGND.n841 8569.5
R975 VGND.n905 VGND.n889 8569.5
R976 VGND.n905 VGND.n904 8569.5
R977 VGND.n839 VGND.n304 8569.5
R978 VGND.n839 VGND.n807 8569.5
R979 VGND.n2606 VGND.n807 8569.5
R980 VGND.n2607 VGND.n2606 8569.5
R981 VGND.n2600 VGND.n293 8569.5
R982 VGND.n2600 VGND.n837 8569.5
R983 VGND.n837 VGND.n836 8569.5
R984 VGND.n836 VGND.n803 8569.5
R985 VGND.n3033 VGND.n279 8569.5
R986 VGND.n799 VGND.n279 8569.5
R987 VGND.n838 VGND.n292 8569.5
R988 VGND.n838 VGND.n794 8569.5
R989 VGND.n2614 VGND.n794 8569.5
R990 VGND.n2614 VGND.n2613 8569.5
R991 VGND.n2632 VGND.n780 7827.71
R992 VGND.n2631 VGND.n780 7827.71
R993 VGND.n3141 VGND.n154 7827.71
R994 VGND.n3141 VGND.n155 7827.71
R995 VGND.n1265 VGND.n1171 7333.74
R996 VGND.n1171 VGND.n1169 7333.74
R997 VGND.n1170 VGND.n1169 7333.74
R998 VGND.n1265 VGND.n1170 7333.74
R999 VGND.n1167 VGND.n1166 7333.74
R1000 VGND.n1168 VGND.n1167 7333.74
R1001 VGND.n1197 VGND.n1168 7333.74
R1002 VGND.n1197 VGND.n1166 7333.74
R1003 VGND.n1196 VGND.n1195 7333.74
R1004 VGND.n1201 VGND.n1196 7333.74
R1005 VGND.n1202 VGND.n1201 7333.74
R1006 VGND.n1202 VGND.n1195 7333.74
R1007 VGND.n165 VGND.n164 7027.48
R1008 VGND.n164 VGND.n160 7027.48
R1009 VGND.n745 VGND.n163 7027.48
R1010 VGND.n745 VGND.n159 7027.48
R1011 VGND.n184 VGND.n178 7027.48
R1012 VGND.n184 VGND.n182 7027.48
R1013 VGND.n755 VGND.n177 7027.48
R1014 VGND.n755 VGND.n181 7027.48
R1015 VGND.n2655 VGND.n760 7027.48
R1016 VGND.n760 VGND.n758 7027.48
R1017 VGND.n765 VGND.n761 7027.48
R1018 VGND.n765 VGND.n764 7027.48
R1019 VGND.n771 VGND.n770 7027.48
R1020 VGND.n771 VGND.n768 7027.48
R1021 VGND.n2620 VGND.n781 7027.48
R1022 VGND.n2630 VGND.n2620 7027.48
R1023 VGND.n193 VGND.n189 7027.48
R1024 VGND.n193 VGND.n187 7027.48
R1025 VGND.n1268 VGND.n1162 6876
R1026 VGND.n1268 VGND.n1267 6876
R1027 VGND.n1267 VGND.n1163 6876
R1028 VGND.n1163 VGND.n1162 6876
R1029 VGND.n1600 VGND.n1599 6384.43
R1030 VGND.n3032 VGND.n195 5693.44
R1031 VGND.n3143 VGND.n3142 5395.46
R1032 VGND.n1465 VGND.n1385 4699.26
R1033 VGND.n1385 VGND.n1383 4699.26
R1034 VGND.n1446 VGND.n1401 4699.26
R1035 VGND.n1447 VGND.n1401 4699.26
R1036 VGND.n1382 VGND.n1380 4699.26
R1037 VGND.n1466 VGND.n1380 4699.26
R1038 VGND.n1440 VGND.n1403 4699.26
R1039 VGND.n1440 VGND.n1402 4699.26
R1040 VGND.n1600 VGND.n1159 4652.5
R1041 VGND.n1965 VGND.n1600 4532.81
R1042 VGND.n153 VGND.n152 4450.15
R1043 VGND.n1421 VGND.n1398 3734.38
R1044 VGND.n1421 VGND.n1393 3734.38
R1045 VGND.n1427 VGND.n1384 3734.38
R1046 VGND.n1427 VGND.n1394 3734.38
R1047 VGND.n1423 VGND.n1418 3734.38
R1048 VGND.n1423 VGND.n1419 3734.38
R1049 VGND.n1429 VGND.n1425 3734.38
R1050 VGND.n1429 VGND.n1379 3734.38
R1051 VGND.n3032 VGND.n3031 3633.95
R1052 VGND.n3106 VGND.n3105 3468.42
R1053 VGND.n3221 VGND.n3220 3382.02
R1054 VGND.n3220 VGND.n3212 3382.02
R1055 VGND.n3213 VGND.n3212 3382.02
R1056 VGND.n3221 VGND.n3213 3382.02
R1057 VGND.n3238 VGND.n50 3382.02
R1058 VGND.n3239 VGND.n50 3382.02
R1059 VGND.n3239 VGND.n49 3382.02
R1060 VGND.n3238 VGND.n49 3382.02
R1061 VGND.n91 VGND.n89 3382.02
R1062 VGND.n3222 VGND.n89 3382.02
R1063 VGND.n3222 VGND.n88 3382.02
R1064 VGND.n91 VGND.n88 3382.02
R1065 VGND.n86 VGND.n47 3382.02
R1066 VGND.n86 VGND.n52 3382.02
R1067 VGND.n3167 VGND.n52 3382.02
R1068 VGND.n3167 VGND.n47 3382.02
R1069 VGND.n3146 VGND.n84 3382.02
R1070 VGND.n3211 VGND.n3146 3382.02
R1071 VGND.n3211 VGND.n3145 3382.02
R1072 VGND.n3145 VGND.n84 3382.02
R1073 VGND.n3175 VGND.n57 3382.02
R1074 VGND.n3175 VGND.n56 3382.02
R1075 VGND.n3165 VGND.n56 3382.02
R1076 VGND.n3165 VGND.n57 3382.02
R1077 VGND.n3148 VGND.n92 3382.02
R1078 VGND.n3148 VGND.n93 3382.02
R1079 VGND.n3156 VGND.n93 3382.02
R1080 VGND.n3156 VGND.n92 3382.02
R1081 VGND.n3155 VGND.n53 3382.02
R1082 VGND.n3155 VGND.n54 3382.02
R1083 VGND.n3187 VGND.n54 3382.02
R1084 VGND.n3187 VGND.n53 3382.02
R1085 VGND.n3106 VGND.n195 3204.72
R1086 VGND.n1568 VGND.n1567 2985.44
R1087 VGND.n100 VGND.n98 2130.64
R1088 VGND.n107 VGND.n100 2130.64
R1089 VGND.n108 VGND.n107 2130.64
R1090 VGND.n108 VGND.n98 2130.64
R1091 VGND.n111 VGND.n94 2130.64
R1092 VGND.n111 VGND.n95 2130.64
R1093 VGND.n116 VGND.n95 2130.64
R1094 VGND.n116 VGND.n94 2130.64
R1095 VGND.n1599 VGND.n1598 1573.32
R1096 VGND.n3265 VGND.n21 1570.81
R1097 VGND.n3265 VGND.n22 1570.81
R1098 VGND.n3262 VGND.n22 1570.81
R1099 VGND.n3262 VGND.n21 1570.81
R1100 VGND.n149 VGND.n118 1570.81
R1101 VGND.n149 VGND.n119 1570.81
R1102 VGND.n144 VGND.n119 1570.81
R1103 VGND.n144 VGND.n118 1570.81
R1104 VGND.n141 VGND.n128 1570.81
R1105 VGND.n130 VGND.n128 1570.81
R1106 VGND.n134 VGND.n130 1570.81
R1107 VGND.n141 VGND.n134 1570.81
R1108 VGND.n132 VGND.n17 1570.81
R1109 VGND.n132 VGND.n18 1570.81
R1110 VGND.n3267 VGND.n18 1570.81
R1111 VGND.n3267 VGND.n17 1570.81
R1112 VGND.n3059 VGND.n238 1133.93
R1113 VGND.n247 VGND.n240 1133.93
R1114 VGND.n3049 VGND.n252 1133.93
R1115 VGND.n264 VGND.n258 1133.93
R1116 VGND.n1143 VGND.n1100 1133.93
R1117 VGND.n1109 VGND.n1101 1133.93
R1118 VGND.n1133 VGND.n1116 1133.93
R1119 VGND.n1127 VGND.n1118 1133.93
R1120 VGND.n258 VGND.n257 1133.93
R1121 VGND.n1118 VGND.n200 1133.93
R1122 VGND.n1133 VGND.n1117 1133.93
R1123 VGND.n1105 VGND.n1101 1133.93
R1124 VGND.n1143 VGND.n208 1133.93
R1125 VGND.n3049 VGND.n256 1133.93
R1126 VGND.n240 VGND.n216 1133.93
R1127 VGND.n3059 VGND.n239 1133.93
R1128 VGND.n3068 VGND.n225 1133.93
R1129 VGND.n3064 VGND.n225 1133.93
R1130 VGND.n238 VGND.n232 1125.27
R1131 VGND.n3054 VGND.n247 1125.27
R1132 VGND.n252 VGND.n248 1125.27
R1133 VGND.n265 VGND.n264 1125.27
R1134 VGND.n1100 VGND.n1093 1125.27
R1135 VGND.n1138 VGND.n1109 1125.27
R1136 VGND.n1116 VGND.n1110 1125.27
R1137 VGND.n1128 VGND.n1127 1125.27
R1138 VGND.n3069 VGND.n3068 1125.27
R1139 VGND.n257 VGND.n209 1118.12
R1140 VGND.n3102 VGND.n200 1118.12
R1141 VGND.n1117 VGND.n201 1118.12
R1142 VGND.n1105 VGND.n207 1118.12
R1143 VGND.n3093 VGND.n208 1118.12
R1144 VGND.n256 VGND.n215 1118.12
R1145 VGND.n3084 VGND.n216 1118.12
R1146 VGND.n239 VGND.n217 1118.12
R1147 VGND.n3064 VGND.n223 1118.12
R1148 VGND.n1598 VGND.t22 1083.1
R1149 VGND.t124 VGND.n1160 1064.96
R1150 VGND.t124 VGND.n1200 1043.41
R1151 VGND.n1446 VGND.n1393 964.88
R1152 VGND.n1452 VGND.n1393 964.88
R1153 VGND.n1452 VGND.n1394 964.88
R1154 VGND.n1394 VGND.n1383 964.88
R1155 VGND.n1447 VGND.n1398 964.88
R1156 VGND.n1451 VGND.n1398 964.88
R1157 VGND.n1451 VGND.n1384 964.88
R1158 VGND.n1465 VGND.n1384 964.88
R1159 VGND.n1419 VGND.n1403 964.88
R1160 VGND.n1419 VGND.n1396 964.88
R1161 VGND.n1396 VGND.n1379 964.88
R1162 VGND.n1466 VGND.n1379 964.88
R1163 VGND.n1418 VGND.n1402 964.88
R1164 VGND.n1418 VGND.n1395 964.88
R1165 VGND.n1425 VGND.n1395 964.88
R1166 VGND.n1425 VGND.n1382 964.88
R1167 VGND.n1582 VGND.n1010 958.264
R1168 VGND.n3079 VGND.n3078 862.23
R1169 VGND.n1472 VGND.n1313 857.529
R1170 VGND.n1474 VGND.n1472 857.529
R1171 VGND.n1474 VGND.n1473 857.529
R1172 VGND.n1473 VGND.n1326 857.529
R1173 VGND.n1373 VGND.n1326 857.529
R1174 VGND.n1373 VGND.n1340 857.529
R1175 VGND.n1482 VGND.n1340 857.529
R1176 VGND.n1484 VGND.n1482 857.529
R1177 VGND.n1484 VGND.n1483 857.529
R1178 VGND.n1483 VGND.n1352 857.529
R1179 VGND.n1369 VGND.n1352 857.529
R1180 VGND.n1493 VGND.n1369 857.529
R1181 VGND.n1493 VGND.n1370 857.529
R1182 VGND.n1370 VGND.n15 857.529
R1183 VGND.n1533 VGND.n1310 857.529
R1184 VGND.n1332 VGND.n1310 857.529
R1185 VGND.n1332 VGND.n1329 857.529
R1186 VGND.n1524 VGND.n1329 857.529
R1187 VGND.n1524 VGND.n1330 857.529
R1188 VGND.n1520 VGND.n1330 857.529
R1189 VGND.n1520 VGND.n1338 857.529
R1190 VGND.n1358 VGND.n1338 857.529
R1191 VGND.n1358 VGND.n1355 857.529
R1192 VGND.n1511 VGND.n1355 857.529
R1193 VGND.n1511 VGND.n1356 857.529
R1194 VGND.n1503 VGND.n1356 857.529
R1195 VGND.n1503 VGND.n1502 857.529
R1196 VGND.n1502 VGND.n1495 857.529
R1197 VGND.n1387 VGND.n1314 857.529
R1198 VGND.n1316 VGND.n1314 857.529
R1199 VGND.n1527 VGND.n1316 857.529
R1200 VGND.n1527 VGND.n1526 857.529
R1201 VGND.n1526 VGND.n1525 857.529
R1202 VGND.n1525 VGND.n1322 857.529
R1203 VGND.n1341 VGND.n1322 857.529
R1204 VGND.n1342 VGND.n1341 857.529
R1205 VGND.n1514 VGND.n1342 857.529
R1206 VGND.n1514 VGND.n1513 857.529
R1207 VGND.n1513 VGND.n1512 857.529
R1208 VGND.n1512 VGND.n1348 857.529
R1209 VGND.n1504 VGND.n1348 857.529
R1210 VGND.n1504 VGND.n1366 857.529
R1211 VGND.n1366 VGND.n1365 857.529
R1212 VGND.n1365 VGND.n14 857.529
R1213 VGND.n3104 VGND.n198 857.529
R1214 VGND.n3100 VGND.n198 857.529
R1215 VGND.n3100 VGND.n3099 857.529
R1216 VGND.n3099 VGND.n3098 857.529
R1217 VGND.n3098 VGND.n203 857.529
R1218 VGND.n3095 VGND.n203 857.529
R1219 VGND.n3095 VGND.n206 857.529
R1220 VGND.n3091 VGND.n206 857.529
R1221 VGND.n3091 VGND.n3090 857.529
R1222 VGND.n3090 VGND.n3089 857.529
R1223 VGND.n3089 VGND.n211 857.529
R1224 VGND.n3086 VGND.n211 857.529
R1225 VGND.n3086 VGND.n214 857.529
R1226 VGND.n3082 VGND.n214 857.529
R1227 VGND.n3082 VGND.n3081 857.529
R1228 VGND.n3081 VGND.n3080 857.529
R1229 VGND.n3080 VGND.n219 857.529
R1230 VGND.n3078 VGND.n219 857.529
R1231 VGND.n1123 VGND.n1089 857.529
R1232 VGND.n1130 VGND.n1123 857.529
R1233 VGND.n1130 VGND.n1111 857.529
R1234 VGND.n1136 VGND.n1111 857.529
R1235 VGND.n1136 VGND.n1104 857.529
R1236 VGND.n1140 VGND.n1104 857.529
R1237 VGND.n1140 VGND.n1094 857.529
R1238 VGND.n1146 VGND.n1094 857.529
R1239 VGND.n1146 VGND.n261 857.529
R1240 VGND.n3046 VGND.n261 857.529
R1241 VGND.n3046 VGND.n249 857.529
R1242 VGND.n3052 VGND.n249 857.529
R1243 VGND.n3052 VGND.n243 857.529
R1244 VGND.n3056 VGND.n243 857.529
R1245 VGND.n3056 VGND.n233 857.529
R1246 VGND.n3062 VGND.n233 857.529
R1247 VGND.n3062 VGND.n230 857.529
R1248 VGND.n3072 VGND.n230 857.529
R1249 VGND.n1120 VGND.n1090 857.529
R1250 VGND.n1121 VGND.n1120 857.529
R1251 VGND.n1131 VGND.n1121 857.529
R1252 VGND.n1131 VGND.n1113 857.529
R1253 VGND.n1135 VGND.n1113 857.529
R1254 VGND.n1135 VGND.n1102 857.529
R1255 VGND.n1141 VGND.n1102 857.529
R1256 VGND.n1141 VGND.n1096 857.529
R1257 VGND.n1145 VGND.n1096 857.529
R1258 VGND.n1145 VGND.n259 857.529
R1259 VGND.n3047 VGND.n259 857.529
R1260 VGND.n3047 VGND.n251 857.529
R1261 VGND.n3051 VGND.n251 857.529
R1262 VGND.n3051 VGND.n241 857.529
R1263 VGND.n3057 VGND.n241 857.529
R1264 VGND.n3057 VGND.n235 857.529
R1265 VGND.n3061 VGND.n235 857.529
R1266 VGND.n3061 VGND.n226 857.529
R1267 VGND.n3073 VGND.n226 857.529
R1268 VGND.n3073 VGND.n227 857.529
R1269 VGND.n1562 VGND.n1276 857.529
R1270 VGND.n1556 VGND.n1276 857.529
R1271 VGND.n1556 VGND.n1288 857.529
R1272 VGND.n1552 VGND.n1288 857.529
R1273 VGND.n1552 VGND.n1291 857.529
R1274 VGND.n1546 VGND.n1291 857.529
R1275 VGND.n1561 VGND.n1279 857.529
R1276 VGND.n1557 VGND.n1279 857.529
R1277 VGND.n1557 VGND.n1284 857.529
R1278 VGND.n1551 VGND.n1284 857.529
R1279 VGND.n1551 VGND.n1295 857.529
R1280 VGND.n1547 VGND.n1295 857.529
R1281 VGND.n2632 VGND.n781 800.225
R1282 VGND.n2628 VGND.n781 800.225
R1283 VGND.n2628 VGND.n770 800.225
R1284 VGND.n2648 VGND.n770 800.225
R1285 VGND.n2648 VGND.n761 800.225
R1286 VGND.n2654 VGND.n761 800.225
R1287 VGND.n2655 VGND.n2654 800.225
R1288 VGND.n2656 VGND.n2655 800.225
R1289 VGND.n2656 VGND.n177 800.225
R1290 VGND.n3120 VGND.n177 800.225
R1291 VGND.n3120 VGND.n178 800.225
R1292 VGND.n3114 VGND.n178 800.225
R1293 VGND.n3114 VGND.n189 800.225
R1294 VGND.n3109 VGND.n189 800.225
R1295 VGND.n3109 VGND.n163 800.225
R1296 VGND.n3135 VGND.n163 800.225
R1297 VGND.n3135 VGND.n165 800.225
R1298 VGND.n165 VGND.n154 800.225
R1299 VGND.n2631 VGND.n2630 800.225
R1300 VGND.n2630 VGND.n2629 800.225
R1301 VGND.n2629 VGND.n768 800.225
R1302 VGND.n2649 VGND.n768 800.225
R1303 VGND.n2649 VGND.n764 800.225
R1304 VGND.n2653 VGND.n764 800.225
R1305 VGND.n2653 VGND.n758 800.225
R1306 VGND.n2657 VGND.n758 800.225
R1307 VGND.n2657 VGND.n181 800.225
R1308 VGND.n3119 VGND.n181 800.225
R1309 VGND.n3119 VGND.n182 800.225
R1310 VGND.n3115 VGND.n182 800.225
R1311 VGND.n3115 VGND.n187 800.225
R1312 VGND.n3108 VGND.n187 800.225
R1313 VGND.n3108 VGND.n159 800.225
R1314 VGND.n3136 VGND.n159 800.225
R1315 VGND.n3136 VGND.n160 800.225
R1316 VGND.n160 VGND.n155 800.225
R1317 VGND.n2651 VGND.n766 791.341
R1318 VGND.n939 VGND.n757 791.341
R1319 VGND.n2659 VGND.n756 791.341
R1320 VGND.n3117 VGND.n185 791.341
R1321 VGND.n746 VGND.n158 791.341
R1322 VGND.n772 VGND.n767 791.341
R1323 VGND.n2624 VGND.n2623 791.341
R1324 VGND.n192 VGND.n186 791.341
R1325 VGND.n3138 VGND.n157 791.341
R1326 VGND.n3111 VGND.n191 787.617
R1327 VGND.n2646 VGND.n2645 787.577
R1328 VGND.n941 VGND.n940 787.577
R1329 VGND.n3122 VGND.n175 787.577
R1330 VGND.n736 VGND.n176 787.577
R1331 VGND.n747 VGND.n166 787.577
R1332 VGND.n774 VGND.n773 787.577
R1333 VGND.n2626 VGND.n2625 787.577
R1334 VGND.n3133 VGND.n3132 787.577
R1335 VGND.n1529 VGND.n1317 776.283
R1336 VGND.n1376 VGND.n1319 776.283
R1337 VGND.n1375 VGND.n1372 776.283
R1338 VGND.n1516 VGND.n1343 776.283
R1339 VGND.n1371 VGND.n1345 776.283
R1340 VGND.n1500 VGND.n1363 776.283
R1341 VGND.n1357 VGND.n1345 776.283
R1342 VGND.n1517 VGND.n1516 776.283
R1343 VGND.n1372 VGND.n1336 776.283
R1344 VGND.n1331 VGND.n1319 776.283
R1345 VGND.n1530 VGND.n1529 776.283
R1346 VGND.n1508 VGND.n1506 776.283
R1347 VGND.n1506 VGND.n1362 776.283
R1348 VGND.n1490 VGND.n1363 776.283
R1349 VGND.n1500 VGND.n1499 774.777
R1350 VGND.n1360 VGND.n1357 774.777
R1351 VGND.n1517 VGND.n1337 774.777
R1352 VGND.n1522 VGND.n1336 774.777
R1353 VGND.n1334 VGND.n1331 774.777
R1354 VGND.n1530 VGND.n1308 774.777
R1355 VGND.n1509 VGND.n1508 774.777
R1356 VGND.n1470 VGND.n1317 765.365
R1357 VGND.n1476 VGND.n1376 765.365
R1358 VGND.n1478 VGND.n1375 765.365
R1359 VGND.n1480 VGND.n1343 765.365
R1360 VGND.n1486 VGND.n1371 765.365
R1361 VGND.n1488 VGND.n1362 765.365
R1362 VGND.n1491 VGND.n1490 765.365
R1363 VGND.n3018 VGND.n292 759.029
R1364 VGND.n3018 VGND.n293 759.029
R1365 VGND.n3016 VGND.n293 759.029
R1366 VGND.n3016 VGND.n304 759.029
R1367 VGND.n304 VGND.n294 759.029
R1368 VGND.n840 VGND.n294 759.029
R1369 VGND.n840 VGND.n303 759.029
R1370 VGND.n842 VGND.n303 759.029
R1371 VGND.n842 VGND.n295 759.029
R1372 VGND.n844 VGND.n295 759.029
R1373 VGND.n844 VGND.n302 759.029
R1374 VGND.n846 VGND.n302 759.029
R1375 VGND.n846 VGND.n296 759.029
R1376 VGND.n848 VGND.n296 759.029
R1377 VGND.n848 VGND.n301 759.029
R1378 VGND.n850 VGND.n301 759.029
R1379 VGND.n850 VGND.n297 759.029
R1380 VGND.n852 VGND.n297 759.029
R1381 VGND.n852 VGND.n300 759.029
R1382 VGND.n854 VGND.n300 759.029
R1383 VGND.n854 VGND.n298 759.029
R1384 VGND.n857 VGND.n788 759.029
R1385 VGND.n944 VGND.n788 759.029
R1386 VGND.n929 VGND.n856 759.029
R1387 VGND.n937 VGND.n856 759.029
R1388 VGND.n938 VGND.n937 759.029
R1389 VGND.n865 VGND.n787 759.029
R1390 VGND.n863 VGND.n787 759.029
R1391 VGND.n863 VGND.n789 759.029
R1392 VGND.n857 VGND.n789 759.029
R1393 VGND.n919 VGND.n864 759.029
R1394 VGND.n927 VGND.n864 759.029
R1395 VGND.n928 VGND.n927 759.029
R1396 VGND.n929 VGND.n928 759.029
R1397 VGND.n872 VGND.n786 759.029
R1398 VGND.n917 VGND.n786 759.029
R1399 VGND.n917 VGND.n790 759.029
R1400 VGND.n865 VGND.n790 759.029
R1401 VGND.n898 VGND.n871 759.029
R1402 VGND.n916 VGND.n871 759.029
R1403 VGND.n920 VGND.n916 759.029
R1404 VGND.n920 VGND.n919 759.029
R1405 VGND.n890 VGND.n785 759.029
R1406 VGND.n896 VGND.n785 759.029
R1407 VGND.n896 VGND.n791 759.029
R1408 VGND.n872 VGND.n791 759.029
R1409 VGND.n904 VGND.n903 759.029
R1410 VGND.n903 VGND.n892 759.029
R1411 VGND.n899 VGND.n892 759.029
R1412 VGND.n899 VGND.n898 759.029
R1413 VGND.n807 VGND.n784 759.029
R1414 VGND.n889 VGND.n784 759.029
R1415 VGND.n889 VGND.n792 759.029
R1416 VGND.n890 VGND.n792 759.029
R1417 VGND.n2608 VGND.n803 759.029
R1418 VGND.n2608 VGND.n2607 759.029
R1419 VGND.n2607 VGND.n806 759.029
R1420 VGND.n904 VGND.n806 759.029
R1421 VGND.n794 VGND.n783 759.029
R1422 VGND.n837 VGND.n783 759.029
R1423 VGND.n837 VGND.n793 759.029
R1424 VGND.n807 VGND.n793 759.029
R1425 VGND.n2618 VGND.n279 759.029
R1426 VGND.n2618 VGND.n794 759.029
R1427 VGND.n292 VGND.n278 759.029
R1428 VGND.n2613 VGND.n802 759.029
R1429 VGND.n2613 VGND.n2612 759.029
R1430 VGND.n2612 VGND.n803 759.029
R1431 VGND.t1 VGND.t107 739.593
R1432 VGND.n1554 VGND.n1289 717.929
R1433 VGND.n1282 VGND.n1274 717.929
R1434 VGND.n1302 VGND.n1296 717.929
R1435 VGND.n1289 VGND.n1283 708.894
R1436 VGND.n1559 VGND.n1282 708.894
R1437 VGND.n1549 VGND.n1296 708.894
R1438 VGND.t91 VGND.n1269 704.476
R1439 VGND.n1537 VGND.n1307 644.495
R1440 VGND.n1537 VGND.n1272 629.587
R1441 VGND.n2852 VGND.n488 601.601
R1442 VGND.n2066 VGND.n397 601.4
R1443 VGND.n398 VGND.n397 600
R1444 VGND.n2852 VGND.n491 599.801
R1445 VGND.n1858 VGND.n1796 585
R1446 VGND.n1864 VGND.n1794 585
R1447 VGND.n1793 VGND.n1783 585
R1448 VGND.n1791 VGND.n1782 585
R1449 VGND.n1874 VGND.n1780 585
R1450 VGND.n1878 VGND.n1771 585
R1451 VGND.n1770 VGND.n1763 585
R1452 VGND.n1768 VGND.n1762 585
R1453 VGND.n1888 VGND.n1760 585
R1454 VGND.n1892 VGND.n1701 585
R1455 VGND.n1751 VGND.n1750 585
R1456 VGND.n1748 VGND.n1747 585
R1457 VGND.n1747 VGND.n1653 585
R1458 VGND.n1753 VGND.n1751 585
R1459 VGND.n1892 VGND.n1891 585
R1460 VGND.n1889 VGND.n1888 585
R1461 VGND.n1762 VGND.n1754 585
R1462 VGND.n1776 VGND.n1763 585
R1463 VGND.n1878 VGND.n1877 585
R1464 VGND.n1875 VGND.n1874 585
R1465 VGND.n1782 VGND.n1777 585
R1466 VGND.n1860 VGND.n1783 585
R1467 VGND.n1864 VGND.n1863 585
R1468 VGND.n1861 VGND.n1858 585
R1469 VGND.n2555 VGND.n2554 585
R1470 VGND.n967 VGND.n715 585
R1471 VGND.n2683 VGND.n715 585
R1472 VGND.n2569 VGND.n961 585
R1473 VGND.n961 VGND.n960 585
R1474 VGND.n2578 VGND.n2577 585
R1475 VGND.n2579 VGND.n2578 585
R1476 VGND.n964 VGND.n962 585
R1477 VGND.n962 VGND.n959 585
R1478 VGND.n2456 VGND.n2454 585
R1479 VGND.n2458 VGND.n2456 585
R1480 VGND.n2559 VGND.n2558 585
R1481 VGND.n2558 VGND.n2557 585
R1482 VGND.n2457 VGND.n2455 585
R1483 VGND.n2556 VGND.n2457 585
R1484 VGND.n2546 VGND.n2481 585
R1485 VGND.n2545 VGND.n2483 585
R1486 VGND.n2545 VGND.n2544 585
R1487 VGND.n2486 VGND.n2482 585
R1488 VGND.n2543 VGND.n2482 585
R1489 VGND.n2541 VGND.n2540 585
R1490 VGND.n2542 VGND.n2541 585
R1491 VGND.n2536 VGND.n2485 585
R1492 VGND.n2485 VGND.n2484 585
R1493 VGND.n2490 VGND.n2488 585
R1494 VGND.n2492 VGND.n2490 585
R1495 VGND.n2531 VGND.n2530 585
R1496 VGND.n2530 VGND.n2529 585
R1497 VGND.n2495 VGND.n2491 585
R1498 VGND.n2528 VGND.n2491 585
R1499 VGND.n2526 VGND.n2525 585
R1500 VGND.n2527 VGND.n2526 585
R1501 VGND.n2522 VGND.n2494 585
R1502 VGND.n2494 VGND.n2493 585
R1503 VGND.n2520 VGND.n2519 585
R1504 VGND.n2519 VGND.n2518 585
R1505 VGND.n2515 VGND.n369 585
R1506 VGND.n371 VGND.n369 585
R1507 VGND.n2934 VGND.n370 585
R1508 VGND.n2934 VGND.n2933 585
R1509 VGND.n665 VGND.n664 585
R1510 VGND.n2957 VGND.n2956 585
R1511 VGND.n2994 VGND.n2993 585
R1512 VGND.n2997 VGND.n319 585
R1513 VGND.n1825 VGND.n1824 585
R1514 VGND.n1830 VGND.n1822 585
R1515 VGND.n1834 VGND.n1819 585
R1516 VGND.n1817 VGND.n1816 585
R1517 VGND.n1840 VGND.n1814 585
R1518 VGND.n1844 VGND.n1808 585
R1519 VGND.n1807 VGND.n1804 585
R1520 VGND.n1850 VGND.n1803 585
R1521 VGND.n1852 VGND.n1802 585
R1522 VGND.n2853 VGND.n490 585
R1523 VGND.n1857 VGND.n388 585
R1524 VGND.n2932 VGND.n388 585
R1525 VGND.n404 VGND.n394 585
R1526 VGND.n405 VGND.n400 585
R1527 VGND.n2920 VGND.n407 585
R1528 VGND.n470 VGND.n408 585
R1529 VGND.n472 VGND.n469 585
R1530 VGND.n2867 VGND.n473 585
R1531 VGND.n2863 VGND.n480 585
R1532 VGND.n482 VGND.n481 585
R1533 VGND.n2858 VGND.n484 585
R1534 VGND.n1797 VGND.n487 585
R1535 VGND.n1856 VGND.n1799 585
R1536 VGND.n1857 VGND.n389 585
R1537 VGND.n2932 VGND.n389 585
R1538 VGND.n1856 VGND.n1855 585
R1539 VGND.n1853 VGND.n1852 585
R1540 VGND.n1850 VGND.n1800 585
R1541 VGND.n1811 VGND.n1804 585
R1542 VGND.n1844 VGND.n1843 585
R1543 VGND.n1841 VGND.n1840 585
R1544 VGND.n1816 VGND.n1812 585
R1545 VGND.n1834 VGND.n1833 585
R1546 VGND.n1831 VGND.n1830 585
R1547 VGND.n1825 VGND.n317 585
R1548 VGND.n2998 VGND.n2997 585
R1549 VGND.n3001 VGND.n3000 585
R1550 VGND.n2939 VGND.n361 585
R1551 VGND.n2940 VGND.n283 585
R1552 VGND.n2943 VGND.n362 585
R1553 VGND.n2944 VGND.n364 585
R1554 VGND.n2948 VGND.n365 585
R1555 VGND.n2950 VGND.n2949 585
R1556 VGND.n663 VGND.n662 585
R1557 VGND.n2935 VGND.n361 585
R1558 VGND.n877 VGND.n876 585
R1559 VGND.n345 VGND.n343 585
R1560 VGND.n2967 VGND.n2966 585
R1561 VGND.n2969 VGND.n342 585
R1562 VGND.n2971 VGND.n2970 585
R1563 VGND.n334 VGND.n332 585
R1564 VGND.n2979 VGND.n2978 585
R1565 VGND.n2981 VGND.n331 585
R1566 VGND.n2983 VGND.n2982 585
R1567 VGND.n324 VGND.n322 585
R1568 VGND.n2990 VGND.n2989 585
R1569 VGND.n2992 VGND.n320 585
R1570 VGND.n355 VGND.n354 585
R1571 VGND.n354 VGND.n283 585
R1572 VGND.n3005 VGND.n3004 585
R1573 VGND.n3008 VGND.n3007 585
R1574 VGND.n312 VGND.n310 585
R1575 VGND.n819 VGND.n306 585
R1576 VGND.n820 VGND.n305 585
R1577 VGND.n823 VGND.n822 585
R1578 VGND.n817 VGND.n812 585
R1579 VGND.n815 VGND.n291 585
R1580 VGND.n814 VGND.n290 585
R1581 VGND.n286 VGND.n284 585
R1582 VGND.n3027 VGND.n3026 585
R1583 VGND.n3029 VGND.n282 585
R1584 VGND.n3003 VGND.n313 585
R1585 VGND.n313 VGND.n283 585
R1586 VGND.n2441 VGND.n2440 585
R1587 VGND.n1575 VGND.n1574 585
R1588 VGND.n1576 VGND.n1575 585
R1589 VGND.n1573 VGND.n997 585
R1590 VGND.n997 VGND.n996 585
R1591 VGND.n2397 VGND.n2396 585
R1592 VGND.n2398 VGND.n2397 585
R1593 VGND.n999 VGND.n995 585
R1594 VGND.n2399 VGND.n995 585
R1595 VGND.n2402 VGND.n2401 585
R1596 VGND.n2401 VGND.n2400 585
R1597 VGND.n2403 VGND.n990 585
R1598 VGND.n990 VGND.n989 585
R1599 VGND.n2412 VGND.n2411 585
R1600 VGND.n2413 VGND.n2412 585
R1601 VGND.n991 VGND.n988 585
R1602 VGND.n2414 VGND.n988 585
R1603 VGND.n2417 VGND.n2416 585
R1604 VGND.n2416 VGND.n2415 585
R1605 VGND.n2418 VGND.n973 585
R1606 VGND.n975 VGND.n973 585
R1607 VGND.n2445 VGND.n2444 585
R1608 VGND.n2444 VGND.n2443 585
R1609 VGND.n974 VGND.n972 585
R1610 VGND.n2442 VGND.n974 585
R1611 VGND.n707 VGND.n703 585
R1612 VGND.n2698 VGND.n2697 585
R1613 VGND.n2697 VGND.n2696 585
R1614 VGND.n706 VGND.n705 585
R1615 VGND.n2695 VGND.n706 585
R1616 VGND.n2693 VGND.n2692 585
R1617 VGND.n2694 VGND.n2693 585
R1618 VGND.n711 VGND.n709 585
R1619 VGND.n709 VGND.n708 585
R1620 VGND.n2686 VGND.n2685 585
R1621 VGND.n2685 VGND.n2684 585
R1622 VGND.n2437 VGND.n2436 585
R1623 VGND.n979 VGND.n977 585
R1624 VGND.n2428 VGND.n984 585
R1625 VGND.n2193 VGND.n2192 585
R1626 VGND.n2196 VGND.n2188 585
R1627 VGND.n2187 VGND.n2185 585
R1628 VGND.n2199 VGND.n693 585
R1629 VGND.n2708 VGND.n2707 585
R1630 VGND.n2710 VGND.n692 585
R1631 VGND.n696 VGND.n692 585
R1632 VGND.n2707 VGND.n2706 585
R1633 VGND.n2199 VGND.n697 585
R1634 VGND.n2185 VGND.n2184 585
R1635 VGND.n2196 VGND.n2195 585
R1636 VGND.n2194 VGND.n2193 585
R1637 VGND.n2428 VGND.n2427 585
R1638 VGND.n979 VGND.n699 585
R1639 VGND.n2704 VGND.n699 585
R1640 VGND.n2436 VGND.n702 585
R1641 VGND.n2025 VGND.n395 585
R1642 VGND.n2033 VGND.n2027 585
R1643 VGND.n2024 VGND.n2021 585
R1644 VGND.n2039 VGND.n2020 585
R1645 VGND.n2043 VGND.n2016 585
R1646 VGND.n2014 VGND.n2012 585
R1647 VGND.n2049 VGND.n2011 585
R1648 VGND.n2053 VGND.n2007 585
R1649 VGND.n2006 VGND.n1069 585
R1650 VGND.n2059 VGND.n1068 585
R1651 VGND.n2063 VGND.n1061 585
R1652 VGND.n1061 VGND.n399 585
R1653 VGND.n2063 VGND.n2062 585
R1654 VGND.n2060 VGND.n2059 585
R1655 VGND.n1069 VGND.n1067 585
R1656 VGND.n2053 VGND.n2052 585
R1657 VGND.n2050 VGND.n2049 585
R1658 VGND.n2017 VGND.n2012 585
R1659 VGND.n2043 VGND.n2042 585
R1660 VGND.n2040 VGND.n2039 585
R1661 VGND.n2021 VGND.n2018 585
R1662 VGND.n2033 VGND.n2032 585
R1663 VGND.n2030 VGND.n395 585
R1664 VGND.n2295 VGND.n2294 585
R1665 VGND.n2293 VGND.n2292 585
R1666 VGND.n2288 VGND.n2078 585
R1667 VGND.n2109 VGND.n2080 585
R1668 VGND.n2111 VGND.n2081 585
R1669 VGND.n2277 VGND.n2112 585
R1670 VGND.n2273 VGND.n2122 585
R1671 VGND.n2126 VGND.n2125 585
R1672 VGND.n2127 VGND.n684 585
R1673 VGND.n2718 VGND.n2717 585
R1674 VGND.n2854 VGND.n2853 585
R1675 VGND.n2856 VGND.n487 585
R1676 VGND.n2858 VGND.n2857 585
R1677 VGND.n481 VGND.n476 585
R1678 VGND.n2864 VGND.n2863 585
R1679 VGND.n2867 VGND.n2866 585
R1680 VGND.n475 VGND.n469 585
R1681 VGND.n408 VGND.n401 585
R1682 VGND.n2921 VGND.n2920 585
R1683 VGND.n2923 VGND.n400 585
R1684 VGND.n2924 VGND.n394 585
R1685 VGND.n488 VGND.n374 585
R1686 VGND.n2786 VGND.n533 585
R1687 VGND.n2792 VGND.n528 585
R1688 VGND.n527 VGND.n522 585
R1689 VGND.n525 VGND.n521 585
R1690 VGND.n2805 VGND.n516 585
R1691 VGND.n2811 VGND.n511 585
R1692 VGND.n510 VGND.n504 585
R1693 VGND.n508 VGND.n503 585
R1694 VGND.n2846 VGND.n499 585
R1695 VGND.n2850 VGND.n494 585
R1696 VGND.n2850 VGND.n2849 585
R1697 VGND.n2847 VGND.n2846 585
R1698 VGND.n2807 VGND.n503 585
R1699 VGND.n2808 VGND.n504 585
R1700 VGND.n2811 VGND.n2810 585
R1701 VGND.n2806 VGND.n2805 585
R1702 VGND.n2788 VGND.n521 585
R1703 VGND.n2789 VGND.n522 585
R1704 VGND.n2792 VGND.n2791 585
R1705 VGND.n2787 VGND.n2786 585
R1706 VGND.n2550 VGND.n2461 585
R1707 VGND.n2460 VGND.n2450 585
R1708 VGND.n2477 VGND.n2463 585
R1709 VGND.n2472 VGND.n2471 585
R1710 VGND.n2757 VGND.n579 585
R1711 VGND.n2749 VGND.n578 585
R1712 VGND.n2752 VGND.n2751 585
R1713 VGND.n2768 VGND.n572 585
R1714 VGND.n2771 VGND.n567 585
R1715 VGND.n2771 VGND.n2770 585
R1716 VGND.n2769 VGND.n2768 585
R1717 VGND.n2753 VGND.n2752 585
R1718 VGND.n2754 VGND.n578 585
R1719 VGND.n2757 VGND.n2756 585
R1720 VGND.n2472 VGND.n581 585
R1721 VGND.n2479 VGND.n2477 585
R1722 VGND.n2480 VGND.n2450 585
R1723 VGND.n2480 VGND.n379 585
R1724 VGND.n2550 VGND.n2549 585
R1725 VGND.n690 VGND.n689 585
R1726 VGND.n2246 VGND.n2217 585
R1727 VGND.n2216 VGND.n2215 585
R1728 VGND.n2239 VGND.n2234 585
R1729 VGND.n2233 VGND.n2232 585
R1730 VGND.n2226 VGND.n2222 585
R1731 VGND.n2221 VGND.n1038 585
R1732 VGND.n2341 VGND.n1035 585
R1733 VGND.n2345 VGND.n1031 585
R1734 VGND.n1027 VGND.n1026 585
R1735 VGND.n2351 VGND.n1025 585
R1736 VGND.n2355 VGND.n1021 585
R1737 VGND.n2711 VGND.n376 585
R1738 VGND.n691 VGND.n376 585
R1739 VGND.n2745 VGND.n2744 585
R1740 VGND.n673 VGND.n588 585
R1741 VGND.n674 VGND.n592 585
R1742 VGND.n2737 VGND.n595 585
R1743 VGND.n2731 VGND.n2730 585
R1744 VGND.n2144 VGND.n603 585
R1745 VGND.n2137 VGND.n2136 585
R1746 VGND.n2140 VGND.n2139 585
R1747 VGND.n2151 VGND.n2141 585
R1748 VGND.n2262 VGND.n679 585
R1749 VGND.n2726 VGND.n2725 585
R1750 VGND.n680 VGND.n678 585
R1751 VGND.n2704 VGND.n698 585
R1752 VGND.n2748 VGND.n582 585
R1753 VGND.n2748 VGND.n2747 585
R1754 VGND.n2960 VGND.n350 585
R1755 VGND.n660 VGND.n659 585
R1756 VGND.n610 VGND.n609 585
R1757 VGND.n612 VGND.n611 585
R1758 VGND.n646 VGND.n616 585
R1759 VGND.n621 VGND.n620 585
R1760 VGND.n637 VGND.n633 585
R1761 VGND.n632 VGND.n631 585
R1762 VGND.n2778 VGND.n544 585
R1763 VGND.n604 VGND.n540 585
R1764 VGND.n2783 VGND.n539 585
R1765 VGND.n538 VGND.n379 585
R1766 VGND.n589 VGND.n374 585
R1767 VGND.n591 VGND.n381 585
R1768 VGND.n2721 VGND.n381 585
R1769 VGND.n2722 VGND.n680 585
R1770 VGND.n2725 VGND.n2724 585
R1771 VGND.n2262 VGND.n682 585
R1772 VGND.n2151 VGND.n2150 585
R1773 VGND.n2148 VGND.n2139 585
R1774 VGND.n2146 VGND.n2137 585
R1775 VGND.n2145 VGND.n2144 585
R1776 VGND.n2731 VGND.n593 585
R1777 VGND.n2738 VGND.n2737 585
R1778 VGND.n2740 VGND.n592 585
R1779 VGND.n2741 VGND.n588 585
R1780 VGND.n2744 VGND.n2743 585
R1781 VGND.n541 VGND.n381 585
R1782 VGND.n2783 VGND.n2782 585
R1783 VGND.n2780 VGND.n540 585
R1784 VGND.n2779 VGND.n2778 585
R1785 VGND.n631 VGND.n622 585
R1786 VGND.n638 VGND.n637 585
R1787 VGND.n640 VGND.n621 585
R1788 VGND.n646 VGND.n645 585
R1789 VGND.n643 VGND.n612 585
R1790 VGND.n642 VGND.n610 585
R1791 VGND.n659 VGND.n352 585
R1792 VGND.n2960 VGND.n2959 585
R1793 VGND.n688 VGND.n381 585
R1794 VGND.n2355 VGND.n2354 585
R1795 VGND.n2352 VGND.n2351 585
R1796 VGND.n1027 VGND.n1024 585
R1797 VGND.n2345 VGND.n2344 585
R1798 VGND.n2342 VGND.n2341 585
R1799 VGND.n2223 VGND.n1038 585
R1800 VGND.n2226 VGND.n2225 585
R1801 VGND.n2232 VGND.n2218 585
R1802 VGND.n2240 VGND.n2239 585
R1803 VGND.n2242 VGND.n2215 585
R1804 VGND.n2246 VGND.n2245 585
R1805 VGND.n2243 VGND.n689 585
R1806 VGND.n2717 VGND.n2716 585
R1807 VGND.n2127 VGND.n687 585
R1808 VGND.n2126 VGND.n2119 585
R1809 VGND.n2274 VGND.n2273 585
R1810 VGND.n2277 VGND.n2276 585
R1811 VGND.n2117 VGND.n2081 585
R1812 VGND.n2080 VGND.n2076 585
R1813 VGND.n2289 VGND.n2288 585
R1814 VGND.n2292 VGND.n2291 585
R1815 VGND.n2295 VGND.n2068 585
R1816 VGND.n2927 VGND.n396 585
R1817 VGND.n399 VGND.n396 585
R1818 VGND.n2927 VGND.n2926 585
R1819 VGND.n2930 VGND.n387 585
R1820 VGND.n2932 VGND.n387 585
R1821 VGND.n2929 VGND.n393 585
R1822 VGND.n2931 VGND.n2930 585
R1823 VGND.n2932 VGND.n2931 585
R1824 VGND.n2929 VGND.n391 585
R1825 VGND.n2873 VGND.n392 585
R1826 VGND.n2882 VGND.n2875 585
R1827 VGND.n2878 VGND.n2877 585
R1828 VGND.n2890 VGND.n460 585
R1829 VGND.n2897 VGND.n456 585
R1830 VGND.n454 VGND.n448 585
R1831 VGND.n453 VGND.n447 585
R1832 VGND.n451 VGND.n450 585
R1833 VGND.n2908 VGND.n439 585
R1834 VGND.n2912 VGND.n433 585
R1835 VGND.n1632 VGND.n1631 585
R1836 VGND.n1935 VGND.n1629 585
R1837 VGND.n1935 VGND.n1934 585
R1838 VGND.n1632 VGND.n435 585
R1839 VGND.n2912 VGND.n2911 585
R1840 VGND.n2909 VGND.n2908 585
R1841 VGND.n450 VGND.n436 585
R1842 VGND.n2893 VGND.n447 585
R1843 VGND.n2894 VGND.n448 585
R1844 VGND.n2897 VGND.n2896 585
R1845 VGND.n2891 VGND.n2890 585
R1846 VGND.n2879 VGND.n2878 585
R1847 VGND.n2882 VGND.n2881 585
R1848 VGND.n392 VGND.n390 585
R1849 VGND.n1628 VGND.n1619 585
R1850 VGND.n1619 VGND.n383 585
R1851 VGND.n1938 VGND.n1937 585
R1852 VGND.n1939 VGND.n1938 585
R1853 VGND.n1620 VGND.n1618 585
R1854 VGND.n1940 VGND.n1618 585
R1855 VGND.n1943 VGND.n1942 585
R1856 VGND.n1942 VGND.n1941 585
R1857 VGND.n1613 VGND.n1610 585
R1858 VGND.n1610 VGND.n1609 585
R1859 VGND.n1950 VGND.n1949 585
R1860 VGND.n1951 VGND.n1950 585
R1861 VGND.n1611 VGND.n1608 585
R1862 VGND.n1952 VGND.n1608 585
R1863 VGND.n1955 VGND.n1954 585
R1864 VGND.n1954 VGND.n1953 585
R1865 VGND.n1604 VGND.n1602 585
R1866 VGND.n1602 VGND.n1601 585
R1867 VGND.n1962 VGND.n1961 585
R1868 VGND.n1963 VGND.n1962 585
R1869 VGND.n1088 VGND.n1084 585
R1870 VGND.n1964 VGND.n1088 585
R1871 VGND.n1967 VGND.n1966 585
R1872 VGND.n1966 VGND.n1965 585
R1873 VGND.n1900 VGND.n1651 585
R1874 VGND.n1904 VGND.n1651 585
R1875 VGND.n1907 VGND.n1906 585
R1876 VGND.n1906 VGND.n1905 585
R1877 VGND.n1649 VGND.n1645 585
R1878 VGND.n1645 VGND.n1644 585
R1879 VGND.n1913 VGND.n1912 585
R1880 VGND.n1914 VGND.n1913 585
R1881 VGND.n1742 VGND.n1642 585
R1882 VGND.n1915 VGND.n1642 585
R1883 VGND.n1918 VGND.n1917 585
R1884 VGND.n1917 VGND.n1916 585
R1885 VGND.n1641 VGND.n1639 585
R1886 VGND.n1643 VGND.n1641 585
R1887 VGND.n1923 VGND.n1635 585
R1888 VGND.n1635 VGND.n1634 585
R1889 VGND.n1927 VGND.n1926 585
R1890 VGND.n1928 VGND.n1927 585
R1891 VGND.n1637 VGND.n1633 585
R1892 VGND.n1929 VGND.n1633 585
R1893 VGND.n1931 VGND.n1627 585
R1894 VGND.n1931 VGND.n1930 585
R1895 VGND.n1932 VGND.n1628 585
R1896 VGND.n1932 VGND.n382 585
R1897 VGND.n3030 VGND.n276 585
R1898 VGND.n3031 VGND.n3030 585
R1899 VGND.n1671 VGND.n281 585
R1900 VGND.n281 VGND.n280 585
R1901 VGND.n1677 VGND.n1676 585
R1902 VGND.n1678 VGND.n1677 585
R1903 VGND.n1668 VGND.n1666 585
R1904 VGND.n1679 VGND.n1666 585
R1905 VGND.n1682 VGND.n1681 585
R1906 VGND.n1681 VGND.n1680 585
R1907 VGND.n1663 VGND.n1660 585
R1908 VGND.n1667 VGND.n1660 585
R1909 VGND.n1691 VGND.n1690 585
R1910 VGND.n1692 VGND.n1691 585
R1911 VGND.n1661 VGND.n1658 585
R1912 VGND.n1693 VGND.n1658 585
R1913 VGND.n1696 VGND.n1695 585
R1914 VGND.n1695 VGND.n1694 585
R1915 VGND.n1655 VGND.n1654 585
R1916 VGND.n1659 VGND.n1654 585
R1917 VGND.n1899 VGND.n1898 585
R1918 VGND.n1899 VGND.n1652 585
R1919 VGND.n1901 VGND.n1900 585
R1920 VGND.n1902 VGND.n1901 585
R1921 VGND.n1020 VGND.n384 585
R1922 VGND.n2357 VGND.n1013 585
R1923 VGND.n2366 VGND.n2365 585
R1924 VGND.n2368 VGND.n1012 585
R1925 VGND.n2371 VGND.n2370 585
R1926 VGND.n2373 VGND.n1006 585
R1927 VGND.n2382 VGND.n2381 585
R1928 VGND.n2384 VGND.n1005 585
R1929 VGND.n2385 VGND.n1001 585
R1930 VGND.n2388 VGND.n2387 585
R1931 VGND.n1003 VGND.n384 585
R1932 VGND.n1572 VGND.n384 585
R1933 VGND.n2318 VGND.n2317 585
R1934 VGND.n2320 VGND.n1060 585
R1935 VGND.n2321 VGND.n1056 585
R1936 VGND.n2324 VGND.n2323 585
R1937 VGND.n1705 VGND.n1058 585
R1938 VGND.n1710 VGND.n1706 585
R1939 VGND.n1730 VGND.n1729 585
R1940 VGND.n1727 VGND.n1726 585
R1941 VGND.n1722 VGND.n1711 585
R1942 VGND.n1717 VGND.n1716 585
R1943 VGND.n1714 VGND.n1016 585
R1944 VGND.n1023 VGND.n384 585
R1945 VGND.n1087 VGND.n384 585
R1946 VGND.n1081 VGND.n1080 585
R1947 VGND.n1976 VGND.n1975 585
R1948 VGND.n1978 VGND.n1077 585
R1949 VGND.n1981 VGND.n1980 585
R1950 VGND.n1074 VGND.n1073 585
R1951 VGND.n1991 VGND.n1990 585
R1952 VGND.n1993 VGND.n1072 585
R1953 VGND.n1999 VGND.n1998 585
R1954 VGND.n1996 VGND.n1064 585
R1955 VGND.n1995 VGND.n1063 585
R1956 VGND.n1066 VGND.n1063 585
R1957 VGND.n3105 VGND.n196 569.73
R1958 VGND.n3097 VGND.n196 569.73
R1959 VGND.n3097 VGND.n3096 569.73
R1960 VGND.n3096 VGND.n205 569.73
R1961 VGND.n3088 VGND.n205 569.73
R1962 VGND.n3088 VGND.n3087 569.73
R1963 VGND.n3087 VGND.n213 569.73
R1964 VGND.n3079 VGND.n221 563.956
R1965 VGND.n1432 VGND.n1430 431.435
R1966 VGND.n1434 VGND.n1424 431.435
R1967 VGND.n1454 VGND.n1391 431.435
R1968 VGND.n1399 VGND.n1392 431.435
R1969 VGND.n1391 VGND.n1386 426.541
R1970 VGND.n1449 VGND.n1399 426.541
R1971 VGND.n1430 VGND.n1378 425.036
R1972 VGND.n1424 VGND.n1417 425.036
R1973 VGND.n3263 VGND.n23 419.183
R1974 VGND.t46 VGND.n51 385.442
R1975 VGND.t46 VGND.n55 385.442
R1976 VGND.t35 VGND.n90 385.442
R1977 VGND.t35 VGND.n3144 385.442
R1978 VGND.n2514 VGND.n2513 352
R1979 VGND.n2673 VGND.n725 347.606
R1980 VGND.t78 VGND.n383 344.533
R1981 VGND.n1904 VGND.n1903 344.533
R1982 VGND.t1 VGND.n2599 340.002
R1983 VGND.t78 VGND.n382 336.834
R1984 VGND.n1903 VGND.n1902 336.834
R1985 VGND.n1903 VGND.n378 336.171
R1986 VGND.n1903 VGND.n377 331.916
R1987 VGND.t78 VGND.n372 164.887
R1988 VGND.t78 VGND.n374 164.887
R1989 VGND.t78 VGND.n376 164.887
R1990 VGND.t78 VGND.n377 327.661
R1991 VGND.n2748 VGND.t78 164.887
R1992 VGND.t78 VGND.n373 164.833
R1993 VGND.t78 VGND.n375 164.833
R1994 VGND.n2704 VGND.t78 164.833
R1995 VGND.t78 VGND.n378 323.404
R1996 VGND.t78 VGND.n379 164.833
R1997 VGND.n2819 VGND.n2818 321.271
R1998 VGND.t22 VGND.n1576 318.815
R1999 VGND.n2951 VGND.n300 307.063
R2000 VGND.n2951 VGND.n298 306.562
R2001 VGND.n2372 VGND.n1010 303.322
R2002 VGND.n1120 VGND.n1119 292.5
R2003 VGND.n1120 VGND.t10 292.5
R2004 VGND.n1132 VGND.n1131 292.5
R2005 VGND.n1131 VGND.t72 292.5
R2006 VGND.n1135 VGND.n1134 292.5
R2007 VGND.t31 VGND.n1135 292.5
R2008 VGND.n1142 VGND.n1141 292.5
R2009 VGND.n1141 VGND.t17 292.5
R2010 VGND.n1145 VGND.n1144 292.5
R2011 VGND.t8 VGND.n1145 292.5
R2012 VGND.n3048 VGND.n3047 292.5
R2013 VGND.n3047 VGND.t16 292.5
R2014 VGND.n3051 VGND.n3050 292.5
R2015 VGND.t12 VGND.n3051 292.5
R2016 VGND.n3058 VGND.n3057 292.5
R2017 VGND.n3057 VGND.t7 292.5
R2018 VGND.n3061 VGND.n3060 292.5
R2019 VGND.t9 VGND.n3061 292.5
R2020 VGND.n3074 VGND.n3073 292.5
R2021 VGND.n3073 VGND.t21 292.5
R2022 VGND.n1091 VGND.n1089 292.5
R2023 VGND.n1089 VGND.t10 292.5
R2024 VGND.n1130 VGND.n1129 292.5
R2025 VGND.t72 VGND.n1130 292.5
R2026 VGND.n1137 VGND.n1136 292.5
R2027 VGND.n1136 VGND.t31 292.5
R2028 VGND.n1140 VGND.n1139 292.5
R2029 VGND.t17 VGND.n1140 292.5
R2030 VGND.n1147 VGND.n1146 292.5
R2031 VGND.n1146 VGND.t8 292.5
R2032 VGND.n3046 VGND.n3045 292.5
R2033 VGND.t16 VGND.n3046 292.5
R2034 VGND.n3053 VGND.n3052 292.5
R2035 VGND.n3052 VGND.t12 292.5
R2036 VGND.n3056 VGND.n3055 292.5
R2037 VGND.t7 VGND.n3056 292.5
R2038 VGND.n3063 VGND.n3062 292.5
R2039 VGND.n3062 VGND.t9 292.5
R2040 VGND.n3072 VGND.n3071 292.5
R2041 VGND.t21 VGND.n3072 292.5
R2042 VGND.n802 VGND.n801 292.5
R2043 VGND.n802 VGND.n188 292.5
R2044 VGND.n2618 VGND.n2617 292.5
R2045 VGND.n2619 VGND.n2618 292.5
R2046 VGND.n795 VGND.n783 292.5
R2047 VGND.n2619 VGND.n783 292.5
R2048 VGND.n2612 VGND.n2611 292.5
R2049 VGND.n2612 VGND.n188 292.5
R2050 VGND.n2609 VGND.n2608 292.5
R2051 VGND.n2608 VGND.n188 292.5
R2052 VGND.n2603 VGND.n793 292.5
R2053 VGND.n2619 VGND.n793 292.5
R2054 VGND.n808 VGND.n784 292.5
R2055 VGND.n2619 VGND.n784 292.5
R2056 VGND.n887 VGND.n806 292.5
R2057 VGND.n806 VGND.n188 292.5
R2058 VGND.n903 VGND.n902 292.5
R2059 VGND.n903 VGND.n188 292.5
R2060 VGND.n908 VGND.n792 292.5
R2061 VGND.n2619 VGND.n792 292.5
R2062 VGND.n910 VGND.n785 292.5
R2063 VGND.n2619 VGND.n785 292.5
R2064 VGND.n900 VGND.n899 292.5
R2065 VGND.n899 VGND.n188 292.5
R2066 VGND.n893 VGND.n871 292.5
R2067 VGND.n871 VGND.n188 292.5
R2068 VGND.n912 VGND.n791 292.5
R2069 VGND.n2619 VGND.n791 292.5
R2070 VGND.n881 VGND.n786 292.5
R2071 VGND.n2619 VGND.n786 292.5
R2072 VGND.n921 VGND.n920 292.5
R2073 VGND.n920 VGND.n188 292.5
R2074 VGND.n923 VGND.n864 292.5
R2075 VGND.n864 VGND.n188 292.5
R2076 VGND.n873 VGND.n790 292.5
R2077 VGND.n2619 VGND.n790 292.5
R2078 VGND.n867 VGND.n787 292.5
R2079 VGND.n2619 VGND.n787 292.5
R2080 VGND.n928 VGND.n860 292.5
R2081 VGND.n928 VGND.n188 292.5
R2082 VGND.n933 VGND.n856 292.5
R2083 VGND.n856 VGND.n188 292.5
R2084 VGND.n861 VGND.n789 292.5
R2085 VGND.n2619 VGND.n789 292.5
R2086 VGND.n858 VGND.n788 292.5
R2087 VGND.n2619 VGND.n788 292.5
R2088 VGND.n938 VGND.n190 292.5
R2089 VGND.n938 VGND.n188 292.5
R2090 VGND.n3017 VGND.n298 292.5
R2091 VGND.n3017 VGND.n300 292.5
R2092 VGND.n367 VGND.n297 292.5
R2093 VGND.n3017 VGND.n297 292.5
R2094 VGND.n874 VGND.n301 292.5
R2095 VGND.n3017 VGND.n301 292.5
R2096 VGND.n2817 VGND.n296 292.5
R2097 VGND.n3017 VGND.n296 292.5
R2098 VGND.n2977 VGND.n302 292.5
R2099 VGND.n3017 VGND.n302 292.5
R2100 VGND.n327 VGND.n295 292.5
R2101 VGND.n3017 VGND.n295 292.5
R2102 VGND.n2995 VGND.n303 292.5
R2103 VGND.n3017 VGND.n303 292.5
R2104 VGND.n311 VGND.n294 292.5
R2105 VGND.n3017 VGND.n294 292.5
R2106 VGND.n3016 VGND.n3015 292.5
R2107 VGND.n3017 VGND.n3016 292.5
R2108 VGND.n3019 VGND.n3018 292.5
R2109 VGND.n3018 VGND.n3017 292.5
R2110 VGND.n285 VGND.n278 292.5
R2111 VGND.n3017 VGND.n278 292.5
R2112 VGND.n3078 VGND.n3077 292.5
R2113 VGND.n3080 VGND.n220 292.5
R2114 VGND.n3080 VGND.n3079 292.5
R2115 VGND.n3083 VGND.n3082 292.5
R2116 VGND.n3082 VGND.n213 292.5
R2117 VGND.n3086 VGND.n3085 292.5
R2118 VGND.n3087 VGND.n3086 292.5
R2119 VGND.n3089 VGND.n212 292.5
R2120 VGND.n3089 VGND.n3088 292.5
R2121 VGND.n3092 VGND.n3091 292.5
R2122 VGND.n3091 VGND.n205 292.5
R2123 VGND.n3095 VGND.n3094 292.5
R2124 VGND.n3096 VGND.n3095 292.5
R2125 VGND.n3098 VGND.n204 292.5
R2126 VGND.n3098 VGND.n3097 292.5
R2127 VGND.n3101 VGND.n3100 292.5
R2128 VGND.n3100 VGND.n196 292.5
R2129 VGND.n3104 VGND.n3103 292.5
R2130 VGND.n3105 VGND.n3104 292.5
R2131 VGND.n1534 VGND.n1533 292.5
R2132 VGND.n1533 VGND.t11 292.5
R2133 VGND.n1333 VGND.n1332 292.5
R2134 VGND.n1332 VGND.t25 292.5
R2135 VGND.n1524 VGND.n1523 292.5
R2136 VGND.t32 VGND.n1524 292.5
R2137 VGND.n1521 VGND.n1520 292.5
R2138 VGND.n1520 VGND.t33 292.5
R2139 VGND.n1359 VGND.n1358 292.5
R2140 VGND.n1358 VGND.t15 292.5
R2141 VGND.n1511 VGND.n1510 292.5
R2142 VGND.t5 VGND.n1511 292.5
R2143 VGND.n1503 VGND.n1361 292.5
R2144 VGND.t45 VGND.n1503 292.5
R2145 VGND.n1498 VGND.n1495 292.5
R2146 VGND.n1495 VGND.t106 292.5
R2147 VGND.n1318 VGND.n1314 292.5
R2148 VGND.t11 VGND.n1314 292.5
R2149 VGND.n1528 VGND.n1527 292.5
R2150 VGND.n1527 VGND.t25 292.5
R2151 VGND.n1525 VGND.n1323 292.5
R2152 VGND.n1525 VGND.t32 292.5
R2153 VGND.n1344 VGND.n1341 292.5
R2154 VGND.t33 VGND.n1341 292.5
R2155 VGND.n1515 VGND.n1514 292.5
R2156 VGND.n1514 VGND.t15 292.5
R2157 VGND.n1512 VGND.n1349 292.5
R2158 VGND.n1512 VGND.t5 292.5
R2159 VGND.n1505 VGND.n1504 292.5
R2160 VGND.n1504 VGND.t45 292.5
R2161 VGND.n1365 VGND.n1364 292.5
R2162 VGND.n1365 VGND.t106 292.5
R2163 VGND.n15 VGND.n13 292.5
R2164 VGND.t106 VGND.n15 292.5
R2165 VGND.n1493 VGND.n1492 292.5
R2166 VGND.t45 VGND.n1493 292.5
R2167 VGND.n1487 VGND.n1352 292.5
R2168 VGND.t5 VGND.n1352 292.5
R2169 VGND.n1485 VGND.n1484 292.5
R2170 VGND.n1484 VGND.t15 292.5
R2171 VGND.n1479 VGND.n1340 292.5
R2172 VGND.t33 VGND.n1340 292.5
R2173 VGND.n1477 VGND.n1326 292.5
R2174 VGND.t32 VGND.n1326 292.5
R2175 VGND.n1475 VGND.n1474 292.5
R2176 VGND.n1474 VGND.t25 292.5
R2177 VGND.n1469 VGND.n1313 292.5
R2178 VGND.t11 VGND.n1313 292.5
R2179 VGND.n1548 VGND.n1547 292.5
R2180 VGND.n1547 VGND.t130 292.5
R2181 VGND.n1551 VGND.n1550 292.5
R2182 VGND.t88 VGND.n1551 292.5
R2183 VGND.n1558 VGND.n1557 292.5
R2184 VGND.n1557 VGND.t99 292.5
R2185 VGND.n1561 VGND.n1560 292.5
R2186 VGND.t20 VGND.n1561 292.5
R2187 VGND.n1563 VGND.n1562 292.5
R2188 VGND.n1562 VGND.t20 292.5
R2189 VGND.n1556 VGND.n1555 292.5
R2190 VGND.t99 VGND.n1556 292.5
R2191 VGND.n1553 VGND.n1552 292.5
R2192 VGND.n1552 VGND.t88 292.5
R2193 VGND.n1546 VGND.n1545 292.5
R2194 VGND.t130 VGND.n1546 292.5
R2195 VGND.n1590 VGND.n1589 285.99
R2196 VGND.n2670 VGND.n2669 283.363
R2197 VGND.n150 VGND.n117 273.339
R2198 VGND.n2714 VGND.n2713 264.301
R2199 VGND.n1994 VGND.n384 264.301
R2200 VGND.n2553 VGND.n2552 264.301
R2201 VGND.n2547 VGND.n2459 264.301
R2202 VGND.n2936 VGND.n283 264.301
R2203 VGND.n2439 VGND.n976 264.301
R2204 VGND.n2700 VGND.n2699 264.301
R2205 VGND.n2720 VGND.n683 264.301
R2206 VGND.n590 VGND.n535 264.301
R2207 VGND.n2784 VGND.n536 264.301
R2208 VGND.n1571 VGND.n1570 264.301
R2209 VGND.n1712 VGND.n1017 264.301
R2210 VGND.n1629 VGND.n1619 259.416
R2211 VGND.n2066 VGND.n396 259.416
R2212 VGND.n691 VGND.n690 259.416
R2213 VGND.n2993 VGND.n2992 259.416
R2214 VGND.n665 VGND.n662 259.416
R2215 VGND.n2747 VGND.n2745 259.416
R2216 VGND.n3030 VGND.n3029 259.416
R2217 VGND.n1748 VGND.n1651 259.416
R2218 VGND.n2854 VGND.n488 259.416
R2219 VGND.n2313 VGND.n1054 258.334
R2220 VGND.n2359 VGND.n1015 258.334
R2221 VGND.n2258 VGND.n2257 258.334
R2222 VGND.n2773 VGND.n547 258.334
R2223 VGND.n1795 VGND.n377 254.34
R2224 VGND.n1792 VGND.n377 254.34
R2225 VGND.n1779 VGND.n377 254.34
R2226 VGND.n1769 VGND.n377 254.34
R2227 VGND.n1759 VGND.n377 254.34
R2228 VGND.n1749 VGND.n377 254.34
R2229 VGND.n1752 VGND.n378 254.34
R2230 VGND.n1890 VGND.n378 254.34
R2231 VGND.n1775 VGND.n378 254.34
R2232 VGND.n1876 VGND.n378 254.34
R2233 VGND.n1859 VGND.n378 254.34
R2234 VGND.n1862 VGND.n378 254.34
R2235 VGND.n2748 VGND.n586 254.34
R2236 VGND.n2548 VGND.n379 254.34
R2237 VGND.n2728 VGND.n666 254.34
R2238 VGND.n2958 VGND.n353 254.34
R2239 VGND.n399 VGND.n321 254.34
R2240 VGND.n1823 VGND.n399 254.34
R2241 VGND.n1818 VGND.n399 254.34
R2242 VGND.n1813 VGND.n399 254.34
R2243 VGND.n1806 VGND.n399 254.34
R2244 VGND.n1801 VGND.n399 254.34
R2245 VGND.n403 VGND.n316 254.34
R2246 VGND.n406 VGND.n316 254.34
R2247 VGND.n471 VGND.n316 254.34
R2248 VGND.n479 VGND.n316 254.34
R2249 VGND.n483 VGND.n316 254.34
R2250 VGND.n1798 VGND.n316 254.34
R2251 VGND.n1854 VGND.n316 254.34
R2252 VGND.n1810 VGND.n316 254.34
R2253 VGND.n1842 VGND.n316 254.34
R2254 VGND.n1832 VGND.n316 254.34
R2255 VGND.n1821 VGND.n316 254.34
R2256 VGND.n2999 VGND.n316 254.34
R2257 VGND.n2937 VGND.n361 254.34
R2258 VGND.n2938 VGND.n283 254.34
R2259 VGND.n2941 VGND.n362 254.34
R2260 VGND.n2942 VGND.n283 254.34
R2261 VGND.n2945 VGND.n283 254.34
R2262 VGND.n2946 VGND.n359 254.34
R2263 VGND.n2947 VGND.n283 254.34
R2264 VGND.n368 VGND.n283 254.34
R2265 VGND.n875 VGND.n283 254.34
R2266 VGND.n2968 VGND.n283 254.34
R2267 VGND.n340 VGND.n283 254.34
R2268 VGND.n2980 VGND.n283 254.34
R2269 VGND.n329 VGND.n283 254.34
R2270 VGND.n2991 VGND.n283 254.34
R2271 VGND.n3006 VGND.n283 254.34
R2272 VGND.n818 VGND.n283 254.34
R2273 VGND.n821 VGND.n283 254.34
R2274 VGND.n816 VGND.n283 254.34
R2275 VGND.n813 VGND.n283 254.34
R2276 VGND.n3028 VGND.n283 254.34
R2277 VGND.n2438 VGND.n376 254.34
R2278 VGND.n2704 VGND.n2701 254.34
R2279 VGND.n983 VGND.n376 254.34
R2280 VGND.n2191 VGND.n376 254.34
R2281 VGND.n2186 VGND.n376 254.34
R2282 VGND.n2709 VGND.n376 254.34
R2283 VGND.n2704 VGND.n2703 254.34
R2284 VGND.n2705 VGND.n2704 254.34
R2285 VGND.n2704 VGND.n701 254.34
R2286 VGND.n2704 VGND.n700 254.34
R2287 VGND.n2026 VGND.n399 254.34
R2288 VGND.n2023 VGND.n399 254.34
R2289 VGND.n2015 VGND.n399 254.34
R2290 VGND.n2010 VGND.n399 254.34
R2291 VGND.n2005 VGND.n399 254.34
R2292 VGND.n2061 VGND.n316 254.34
R2293 VGND.n2051 VGND.n316 254.34
R2294 VGND.n2009 VGND.n316 254.34
R2295 VGND.n2041 VGND.n316 254.34
R2296 VGND.n2031 VGND.n316 254.34
R2297 VGND.n2029 VGND.n316 254.34
R2298 VGND.n2070 VGND.n373 254.34
R2299 VGND.n2071 VGND.n373 254.34
R2300 VGND.n2110 VGND.n373 254.34
R2301 VGND.n2121 VGND.n373 254.34
R2302 VGND.n2124 VGND.n373 254.34
R2303 VGND.n2719 VGND.n373 254.34
R2304 VGND.n2855 VGND.n399 254.34
R2305 VGND.n486 VGND.n399 254.34
R2306 VGND.n2865 VGND.n399 254.34
R2307 VGND.n474 VGND.n399 254.34
R2308 VGND.n2922 VGND.n399 254.34
R2309 VGND.n2925 VGND.n399 254.34
R2310 VGND.n2848 VGND.n375 254.34
R2311 VGND.n532 VGND.n374 254.34
R2312 VGND.n526 VGND.n374 254.34
R2313 VGND.n515 VGND.n374 254.34
R2314 VGND.n509 VGND.n374 254.34
R2315 VGND.n498 VGND.n374 254.34
R2316 VGND.n496 VGND.n375 254.34
R2317 VGND.n2809 VGND.n375 254.34
R2318 VGND.n513 VGND.n375 254.34
R2319 VGND.n2790 VGND.n375 254.34
R2320 VGND.n530 VGND.n375 254.34
R2321 VGND.n2748 VGND.n585 254.34
R2322 VGND.n2748 VGND.n584 254.34
R2323 VGND.n2750 VGND.n2748 254.34
R2324 VGND.n2748 VGND.n583 254.34
R2325 VGND.n569 VGND.n379 254.34
R2326 VGND.n570 VGND.n379 254.34
R2327 VGND.n2755 VGND.n379 254.34
R2328 VGND.n2478 VGND.n379 254.34
R2329 VGND.n2728 VGND.n667 254.34
R2330 VGND.n2728 VGND.n668 254.34
R2331 VGND.n2728 VGND.n669 254.34
R2332 VGND.n2728 VGND.n670 254.34
R2333 VGND.n2728 VGND.n671 254.34
R2334 VGND.n2728 VGND.n672 254.34
R2335 VGND.n2713 VGND.n2712 254.34
R2336 VGND.n2728 VGND.n587 254.34
R2337 VGND.n2728 VGND.n675 254.34
R2338 VGND.n2729 VGND.n2728 254.34
R2339 VGND.n2728 VGND.n676 254.34
R2340 VGND.n2728 VGND.n677 254.34
R2341 VGND.n2728 VGND.n2727 254.34
R2342 VGND.n2702 VGND.n683 254.34
R2343 VGND.n2746 VGND.n535 254.34
R2344 VGND.n2728 VGND.n661 254.34
R2345 VGND.n2728 VGND.n608 254.34
R2346 VGND.n2728 VGND.n607 254.34
R2347 VGND.n2728 VGND.n606 254.34
R2348 VGND.n2728 VGND.n605 254.34
R2349 VGND.n2784 VGND.n537 254.34
R2350 VGND.n2723 VGND.n353 254.34
R2351 VGND.n2149 VGND.n353 254.34
R2352 VGND.n2147 VGND.n353 254.34
R2353 VGND.n2142 VGND.n353 254.34
R2354 VGND.n2739 VGND.n353 254.34
R2355 VGND.n2742 VGND.n353 254.34
R2356 VGND.n2781 VGND.n353 254.34
R2357 VGND.n542 VGND.n353 254.34
R2358 VGND.n639 VGND.n353 254.34
R2359 VGND.n644 VGND.n353 254.34
R2360 VGND.n641 VGND.n353 254.34
R2361 VGND.n2353 VGND.n353 254.34
R2362 VGND.n2343 VGND.n353 254.34
R2363 VGND.n1033 VGND.n353 254.34
R2364 VGND.n2224 VGND.n353 254.34
R2365 VGND.n2241 VGND.n353 254.34
R2366 VGND.n2244 VGND.n353 254.34
R2367 VGND.n2715 VGND.n372 254.34
R2368 VGND.n2118 VGND.n372 254.34
R2369 VGND.n2275 VGND.n372 254.34
R2370 VGND.n2116 VGND.n372 254.34
R2371 VGND.n2290 VGND.n372 254.34
R2372 VGND.n2067 VGND.n372 254.34
R2373 VGND.n2874 VGND.n385 254.34
R2374 VGND.n2876 VGND.n385 254.34
R2375 VGND.n455 VGND.n385 254.34
R2376 VGND.n452 VGND.n385 254.34
R2377 VGND.n438 VGND.n385 254.34
R2378 VGND.n1630 VGND.n385 254.34
R2379 VGND.n1933 VGND.n386 254.34
R2380 VGND.n2910 VGND.n386 254.34
R2381 VGND.n2892 VGND.n386 254.34
R2382 VGND.n2895 VGND.n386 254.34
R2383 VGND.n458 VGND.n386 254.34
R2384 VGND.n2880 VGND.n386 254.34
R2385 VGND.n1019 VGND.n1017 254.34
R2386 VGND.n1018 VGND.n384 254.34
R2387 VGND.n2367 VGND.n384 254.34
R2388 VGND.n2369 VGND.n384 254.34
R2389 VGND.n2383 VGND.n384 254.34
R2390 VGND.n2386 VGND.n384 254.34
R2391 VGND.n2319 VGND.n384 254.34
R2392 VGND.n2322 VGND.n384 254.34
R2393 VGND.n1709 VGND.n384 254.34
R2394 VGND.n1728 VGND.n384 254.34
R2395 VGND.n1715 VGND.n384 254.34
R2396 VGND.n1713 VGND.n384 254.34
R2397 VGND.n1086 VGND.n1083 254.34
R2398 VGND.n1085 VGND.n384 254.34
R2399 VGND.n1977 VGND.n384 254.34
R2400 VGND.n1979 VGND.n384 254.34
R2401 VGND.n1992 VGND.n384 254.34
R2402 VGND.n1997 VGND.n384 254.34
R2403 VGND.n2675 VGND.n2674 252.327
R2404 VGND.n2508 VGND.n2507 250
R2405 VGND.n2987 VGND.n325 250
R2406 VGND.n1966 VGND.n1087 249.663
R2407 VGND.n2318 VGND.n1061 249.663
R2408 VGND.n1021 VGND.n1020 249.663
R2409 VGND.n491 VGND.n490 249.663
R2410 VGND.n539 VGND.n538 249.663
R2411 VGND.n698 VGND.n678 249.663
R2412 VGND.n1901 VGND.n1653 249.663
R2413 VGND.n1934 VGND.n1932 249.663
R2414 VGND.n2926 VGND.n398 249.663
R2415 VGND.n171 VGND.t29 232.444
R2416 VGND.n1083 VGND.n1079 223.341
R2417 VGND.n2883 VGND.n425 221.667
R2418 VGND.n1866 VGND.n1786 221.667
R2419 VGND.n624 VGND.n623 221.667
R2420 VGND.n2057 VGND.n2003 221.667
R2421 VGND.n2265 VGND.n2264 221.667
R2422 VGND.n1707 VGND.n1009 218.376
R2423 VGND.n1079 VGND.n1078 204.412
R2424 VGND.n99 VGND.n51 204.088
R2425 VGND.n2372 VGND.n1009 204.024
R2426 VGND.n2818 VGND.n351 199.315
R2427 VGND.n1203 VGND.n1190 197.969
R2428 VGND.n393 VGND.n387 197
R2429 VGND.n2440 VGND.n974 197
R2430 VGND.n2957 VGND.n354 197
R2431 VGND.n2935 VGND.n2934 197
R2432 VGND.n2554 VGND.n2457 197
R2433 VGND.n3000 VGND.n313 197
R2434 VGND.n1799 VGND.n388 197
R2435 VGND.n2743 VGND.n591 197
R2436 VGND.n2243 VGND.n688 197
R2437 VGND.n2951 VGND.n363 196.268
R2438 VGND.n2951 VGND.n366 196.268
R2439 VGND.n117 VGND.t42 193.48
R2440 VGND.n110 VGND.t42 193.48
R2441 VGND.n109 VGND.t118 193.48
R2442 VGND.n99 VGND.t118 193.48
R2443 VGND.n2062 VGND.n1066 187.249
R2444 VGND.n1575 VGND.n1572 187.249
R2445 VGND.n2782 VGND.n541 187.249
R2446 VGND.n2546 VGND.n2545 187.249
R2447 VGND.n2697 VGND.n703 187.249
R2448 VGND.n1855 VGND.n389 187.249
R2449 VGND.n2931 VGND.n391 187.249
R2450 VGND.n2722 VGND.n2721 187.249
R2451 VGND.n2354 VGND.n1023 187.249
R2452 VGND.n2728 VGND.n353 185.6
R2453 VGND.n399 VGND.n316 185.6
R2454 VGND.n1707 VGND.n1062 185.018
R2455 VGND.n1788 VGND.n485 185
R2456 VGND.n2860 VGND.n2859 185
R2457 VGND.n2862 VGND.n2861 185
R2458 VGND.n478 VGND.n477 185
R2459 VGND.n2868 VGND.n411 185
R2460 VGND.n2917 VGND.n410 185
R2461 VGND.n2919 VGND.n2918 185
R2462 VGND.n423 VGND.n402 185
R2463 VGND.n425 VGND.n424 185
R2464 VGND.t84 VGND.n425 185
R2465 VGND.n1675 VGND.n1674 185
R2466 VGND.n1673 VGND.n1669 185
R2467 VGND.n1673 VGND.t82 185
R2468 VGND.n1672 VGND.n1665 185
R2469 VGND.n1684 VGND.n1683 185
R2470 VGND.n1689 VGND.n1688 185
R2471 VGND.n1686 VGND.n1662 185
R2472 VGND.n1685 VGND.n1657 185
R2473 VGND.n1698 VGND.n1697 185
R2474 VGND.n1897 VGND.n1896 185
R2475 VGND.n1909 VGND.n1908 185
R2476 VGND.n1911 VGND.n1910 185
R2477 VGND.n1648 VGND.n1647 185
R2478 VGND.n1646 VGND.n1640 185
R2479 VGND.n1920 VGND.n1919 185
R2480 VGND.n1922 VGND.n1921 185
R2481 VGND.n1925 VGND.n1924 185
R2482 VGND.n1638 VGND.n422 185
R2483 VGND.t84 VGND.n422 185
R2484 VGND.n1636 VGND.n430 185
R2485 VGND.n1790 VGND.n1789 185
R2486 VGND.n1871 VGND.n1870 185
R2487 VGND.n1873 VGND.n1872 185
R2488 VGND.n1774 VGND.n1773 185
R2489 VGND.n1772 VGND.n1767 185
R2490 VGND.n1885 VGND.n1884 185
R2491 VGND.n1887 VGND.n1886 185
R2492 VGND.n1757 VGND.n1756 185
R2493 VGND.n1755 VGND.n1700 185
R2494 VGND.n1894 VGND.n1893 185
R2495 VGND.n1758 VGND.n1699 185
R2496 VGND.n1765 VGND.n1761 185
R2497 VGND.n1883 VGND.n1882 185
R2498 VGND.n1880 VGND.n1879 185
R2499 VGND.n1778 VGND.n1766 185
R2500 VGND.n1785 VGND.n1781 185
R2501 VGND.n1869 VGND.n1868 185
R2502 VGND.n1866 VGND.n1865 185
R2503 VGND.n318 VGND.n309 185
R2504 VGND.n1829 VGND.n1828 185
R2505 VGND.n1826 VGND.n1820 185
R2506 VGND.n1836 VGND.n1835 185
R2507 VGND.n1839 VGND.n1838 185
R2508 VGND.n1809 VGND.n1805 185
R2509 VGND.n1846 VGND.n1845 185
R2510 VGND.n1846 VGND.t82 185
R2511 VGND.n1849 VGND.n1848 185
R2512 VGND.n1851 VGND.n1786 185
R2513 VGND.n3010 VGND.n3009 185
R2514 VGND.n3012 VGND.n308 185
R2515 VGND.n3014 VGND.n3013 185
R2516 VGND.n826 VGND.n825 185
R2517 VGND.n828 VGND.n827 185
R2518 VGND.n811 VGND.n289 185
R2519 VGND.n3021 VGND.n3020 185
R2520 VGND.n3023 VGND.n288 185
R2521 VGND.n3025 VGND.n3024 185
R2522 VGND.n2509 VGND.n2508 185
R2523 VGND.n2965 VGND.n2964 185
R2524 VGND.n347 VGND.n344 185
R2525 VGND.n341 VGND.n338 185
R2526 VGND.n2973 VGND.n2972 185
R2527 VGND.n2976 VGND.n2975 185
R2528 VGND.n337 VGND.n336 185
R2529 VGND.n330 VGND.n326 185
R2530 VGND.n2985 VGND.n2984 185
R2531 VGND.n2988 VGND.n2987 185
R2532 VGND.n2819 VGND.n325 185
R2533 VGND.t85 VGND.n325 185
R2534 VGND.n2822 VGND.n2821 185
R2535 VGND.n2823 VGND.n2816 185
R2536 VGND.n2825 VGND.n2824 185
R2537 VGND.n2827 VGND.n2815 185
R2538 VGND.n2830 VGND.n2829 185
R2539 VGND.n2831 VGND.n2814 185
R2540 VGND.n2833 VGND.n2832 185
R2541 VGND.n2833 VGND.t85 185
R2542 VGND.n2834 VGND.n492 185
R2543 VGND.n2562 VGND.n2560 185
R2544 VGND.n2453 VGND.n965 185
R2545 VGND.n2576 VGND.n2575 185
R2546 VGND.n2573 VGND.n963 185
R2547 VGND.n2572 VGND.n2570 185
R2548 VGND.n714 VGND.n713 185
R2549 VGND.n2517 VGND.n2516 185
R2550 VGND.n2521 VGND.n555 185
R2551 VGND.t79 VGND.n555 185
R2552 VGND.n2524 VGND.n2523 185
R2553 VGND.n2498 VGND.n2497 185
R2554 VGND.n2496 VGND.n2489 185
R2555 VGND.n2533 VGND.n2532 185
R2556 VGND.n2535 VGND.n2534 185
R2557 VGND.n2539 VGND.n2538 185
R2558 VGND.n2537 VGND.n2487 185
R2559 VGND.n2359 VGND.n2358 185
R2560 VGND.n2361 VGND.n1014 185
R2561 VGND.n2364 VGND.n2363 185
R2562 VGND.n1011 VGND.n1008 185
R2563 VGND.n2375 VGND.n2374 185
R2564 VGND.n2377 VGND.n1007 185
R2565 VGND.n2380 VGND.n2379 185
R2566 VGND.n1004 VGND.n1000 185
R2567 VGND.n2390 VGND.n2389 185
R2568 VGND.n2422 VGND.n971 185
R2569 VGND.n2420 VGND.n2419 185
R2570 VGND.n987 VGND.n986 185
R2571 VGND.n2410 VGND.n2409 185
R2572 VGND.n2407 VGND.n992 185
R2573 VGND.n2405 VGND.n2404 185
R2574 VGND.n994 VGND.n993 185
R2575 VGND.n2395 VGND.n2394 185
R2576 VGND.n2392 VGND.n998 185
R2577 VGND.n2688 VGND.n2687 185
R2578 VGND.n2691 VGND.n2690 185
R2579 VGND.n712 VGND.n710 185
R2580 VGND.n2423 VGND.n978 185
R2581 VGND.n2426 VGND.n2425 185
R2582 VGND.n985 VGND.n982 185
R2583 VGND.n2189 VGND.n2183 185
R2584 VGND.n2208 VGND.n2207 185
R2585 VGND.n2210 VGND.n2181 185
R2586 VGND.n2211 VGND.n695 185
R2587 VGND.n2213 VGND.n2180 185
R2588 VGND.n2255 VGND.n2254 185
R2589 VGND.n2257 VGND.n2256 185
R2590 VGND.n2198 VGND.n694 185
R2591 VGND.n2201 VGND.n2200 185
R2592 VGND.n2203 VGND.n2197 185
R2593 VGND.n2206 VGND.n2205 185
R2594 VGND.n2190 VGND.n981 185
R2595 VGND.n2430 VGND.n2429 185
R2596 VGND.n2432 VGND.n980 185
R2597 VGND.n2435 VGND.n2434 185
R2598 VGND.n1626 VGND.n1625 185
R2599 VGND.n1617 VGND.n1616 185
R2600 VGND.n1616 VGND.t81 185
R2601 VGND.n1945 VGND.n1944 185
R2602 VGND.n1948 VGND.n1947 185
R2603 VGND.n1615 VGND.n1612 185
R2604 VGND.n1607 VGND.n1606 185
R2605 VGND.n1957 VGND.n1956 185
R2606 VGND.n1960 VGND.n1959 185
R2607 VGND.n1605 VGND.n1603 185
R2608 VGND.n1970 VGND.n1969 185
R2609 VGND.n1973 VGND.n1972 185
R2610 VGND.n1974 VGND.n1076 185
R2611 VGND.n1983 VGND.n1982 185
R2612 VGND.n1985 VGND.n1075 185
R2613 VGND.n1988 VGND.n1987 185
R2614 VGND.n1989 VGND.n1071 185
R2615 VGND.n2001 VGND.n2000 185
R2616 VGND.n2003 VGND.n1070 185
R2617 VGND.n2028 VGND.n466 185
R2618 VGND.n2035 VGND.n2034 185
R2619 VGND.n2038 VGND.n2037 185
R2620 VGND.n2019 VGND.n2013 185
R2621 VGND.n2045 VGND.n2044 185
R2622 VGND.n2048 VGND.n2047 185
R2623 VGND.n2008 VGND.n2004 185
R2624 VGND.n2004 VGND.t81 185
R2625 VGND.n2055 VGND.n2054 185
R2626 VGND.n2058 VGND.n2057 185
R2627 VGND.n1059 VGND.n1054 185
R2628 VGND.n2326 VGND.n2325 185
R2629 VGND.n1057 VGND.n1055 185
R2630 VGND.n1734 VGND.n1733 185
R2631 VGND.n1732 VGND.n1731 185
R2632 VGND.n1723 VGND.n1708 185
R2633 VGND.n1725 VGND.n1724 185
R2634 VGND.n1721 VGND.n1720 185
R2635 VGND.n1719 VGND.n1718 185
R2636 VGND.n2086 VGND.n493 185
R2637 VGND.n2089 VGND.n2088 185
R2638 VGND.n2090 VGND.n2084 185
R2639 VGND.n2092 VGND.n2091 185
R2640 VGND.n2094 VGND.n2083 185
R2641 VGND.n2097 VGND.n2096 185
R2642 VGND.n2098 VGND.n2082 185
R2643 VGND.n2100 VGND.n2099 185
R2644 VGND.n2100 VGND.t77 185
R2645 VGND.n2101 VGND.n2065 185
R2646 VGND.n2298 VGND.n2297 185
R2647 VGND.n2300 VGND.n2299 185
R2648 VGND.n2302 VGND.n2301 185
R2649 VGND.n2304 VGND.n2303 185
R2650 VGND.n2306 VGND.n2305 185
R2651 VGND.n2308 VGND.n2307 185
R2652 VGND.n2310 VGND.n2309 185
R2653 VGND.n2312 VGND.n2311 185
R2654 VGND.n2314 VGND.n2313 185
R2655 VGND.n2248 VGND.n2247 185
R2656 VGND.n2270 VGND.n2269 185
R2657 VGND.n2272 VGND.n2271 185
R2658 VGND.n2115 VGND.n2114 185
R2659 VGND.n2113 VGND.n2108 185
R2660 VGND.n2285 VGND.n2284 185
R2661 VGND.n2287 VGND.n2286 185
R2662 VGND.n2075 VGND.n2074 185
R2663 VGND.n2073 VGND.n2069 185
R2664 VGND.n2103 VGND.n2072 185
R2665 VGND.n2104 VGND.n2077 185
R2666 VGND.n2106 VGND.n2079 185
R2667 VGND.n2282 VGND.n2281 185
R2668 VGND.n2279 VGND.n2278 185
R2669 VGND.n2120 VGND.n2107 185
R2670 VGND.n2129 VGND.n2123 185
R2671 VGND.n2268 VGND.n2267 185
R2672 VGND.n2265 VGND.n685 185
R2673 VGND.n2157 VGND.n529 185
R2674 VGND.n524 VGND.n520 185
R2675 VGND.n2801 VGND.n2800 185
R2676 VGND.n2804 VGND.n2803 185
R2677 VGND.n519 VGND.n512 185
R2678 VGND.n506 VGND.n502 185
R2679 VGND.n2842 VGND.n2841 185
R2680 VGND.n2845 VGND.n2844 185
R2681 VGND.n501 VGND.n495 185
R2682 VGND.n2836 VGND.n497 185
R2683 VGND.n2837 VGND.n500 185
R2684 VGND.n2840 VGND.n2839 185
R2685 VGND.n2813 VGND.n2812 185
R2686 VGND.n2795 VGND.n514 185
R2687 VGND.n2796 VGND.n517 185
R2688 VGND.n2799 VGND.n2798 185
R2689 VGND.n2794 VGND.n2793 185
R2690 VGND.n623 VGND.n531 185
R2691 VGND.n2564 VGND.n2563 185
R2692 VGND.n2476 VGND.n2475 185
R2693 VGND.n2474 VGND.n2473 185
R2694 VGND.n580 VGND.n577 185
R2695 VGND.n2763 VGND.n2762 185
R2696 VGND.n2765 VGND.n576 185
R2697 VGND.n2767 VGND.n2766 185
R2698 VGND.n597 VGND.n568 185
R2699 VGND.n598 VGND.n566 185
R2700 VGND.n2773 VGND.n2772 185
R2701 VGND.n571 VGND.n565 185
R2702 VGND.n574 VGND.n573 185
R2703 VGND.n2759 VGND.n2758 185
R2704 VGND.n2761 VGND.n2760 185
R2705 VGND.n2470 VGND.n2469 185
R2706 VGND.n2468 VGND.n2462 185
R2707 VGND.n2466 VGND.n2465 185
R2708 VGND.n2464 VGND.n2451 185
R2709 VGND.n2252 VGND.n2251 185
R2710 VGND.n2238 VGND.n2214 185
R2711 VGND.n2231 VGND.n2230 185
R2712 VGND.n2228 VGND.n2227 185
R2713 VGND.n2334 VGND.n2333 185
R2714 VGND.n2340 VGND.n2339 185
R2715 VGND.n2337 VGND.n1032 185
R2716 VGND.n2336 VGND.n1030 185
R2717 VGND.n2350 VGND.n1015 185
R2718 VGND.n2158 VGND.n600 185
R2719 VGND.n2736 VGND.n2735 185
R2720 VGND.n2733 VGND.n2732 185
R2721 VGND.n2143 VGND.n601 185
R2722 VGND.n2175 VGND.n2174 185
R2723 VGND.n2172 VGND.n2170 185
R2724 VGND.n2152 VGND.n2132 185
R2725 VGND.n2261 VGND.n2260 185
R2726 VGND.n2258 VGND.n681 185
R2727 VGND.n2507 VGND.n349 185
R2728 VGND.n657 VGND.n656 185
R2729 VGND.n655 VGND.n654 185
R2730 VGND.n619 VGND.n618 185
R2731 VGND.n617 VGND.n615 185
R2732 VGND.n636 VGND.n635 185
R2733 VGND.n630 VGND.n548 185
R2734 VGND.n2777 VGND.n2776 185
R2735 VGND.n547 VGND.n546 185
R2736 VGND.t79 VGND.n547 185
R2737 VGND.n2250 VGND.n2249 185
R2738 VGND.n2237 VGND.n2236 185
R2739 VGND.n2235 VGND.n2219 185
R2740 VGND.n2220 VGND.n1039 185
R2741 VGND.n2332 VGND.n2331 185
R2742 VGND.n2329 VGND.n1036 185
R2743 VGND.n2328 VGND.n1034 185
R2744 VGND.n2347 VGND.n2346 185
R2745 VGND.n2349 VGND.n2348 185
R2746 VGND.n2160 VGND.n2159 185
R2747 VGND.n2162 VGND.n596 185
R2748 VGND.n2163 VGND.n594 185
R2749 VGND.n2165 VGND.n602 185
R2750 VGND.n2166 VGND.n2138 185
R2751 VGND.n2169 VGND.n2168 185
R2752 VGND.n2155 VGND.n2153 185
R2753 VGND.n2131 VGND.n2130 185
R2754 VGND.n2264 VGND.n2263 185
R2755 VGND.n2264 VGND.t77 185
R2756 VGND.n2962 VGND.n2961 185
R2757 VGND.n658 VGND.n348 185
R2758 VGND.n653 VGND.n652 185
R2759 VGND.n650 VGND.n613 185
R2760 VGND.n648 VGND.n647 185
R2761 VGND.n634 VGND.n614 185
R2762 VGND.n629 VGND.n628 185
R2763 VGND.n626 VGND.n545 185
R2764 VGND.n624 VGND.n543 185
R2765 VGND.n2886 VGND.n2885 185
R2766 VGND.n2889 VGND.n2888 185
R2767 VGND.n465 VGND.n457 185
R2768 VGND.n449 VGND.n443 185
R2769 VGND.n2903 VGND.n2902 185
R2770 VGND.n2905 VGND.n442 185
R2771 VGND.n2907 VGND.n2906 185
R2772 VGND.n1622 VGND.n1621 185
R2773 VGND.n1623 VGND.n432 185
R2774 VGND.n2914 VGND.n2913 185
R2775 VGND.n437 VGND.n431 185
R2776 VGND.n444 VGND.n440 185
R2777 VGND.n446 VGND.n445 185
R2778 VGND.n2901 VGND.n2900 185
R2779 VGND.n2899 VGND.n2898 185
R2780 VGND.n461 VGND.n459 185
R2781 VGND.n463 VGND.n462 185
R2782 VGND.n2884 VGND.n2883 185
R2783 VGND.n1976 VGND.n1080 175.546
R2784 VGND.n1980 VGND.n1978 175.546
R2785 VGND.n1991 VGND.n1073 175.546
R2786 VGND.n1998 VGND.n1993 175.546
R2787 VGND.n1996 VGND.n1995 175.546
R2788 VGND.n1966 VGND.n1088 175.546
R2789 VGND.n1962 VGND.n1088 175.546
R2790 VGND.n1962 VGND.n1602 175.546
R2791 VGND.n1954 VGND.n1602 175.546
R2792 VGND.n1954 VGND.n1608 175.546
R2793 VGND.n1950 VGND.n1608 175.546
R2794 VGND.n1950 VGND.n1610 175.546
R2795 VGND.n1942 VGND.n1610 175.546
R2796 VGND.n1942 VGND.n1618 175.546
R2797 VGND.n1938 VGND.n1618 175.546
R2798 VGND.n1938 VGND.n1619 175.546
R2799 VGND.n1631 VGND.n433 175.546
R2800 VGND.n451 VGND.n439 175.546
R2801 VGND.n454 VGND.n453 175.546
R2802 VGND.n460 VGND.n456 175.546
R2803 VGND.n2877 VGND.n2875 175.546
R2804 VGND.n2060 VGND.n1067 175.546
R2805 VGND.n2052 VGND.n2050 175.546
R2806 VGND.n2042 VGND.n2017 175.546
R2807 VGND.n2040 VGND.n2018 175.546
R2808 VGND.n2032 VGND.n2030 175.546
R2809 VGND.n2321 VGND.n2320 175.546
R2810 VGND.n2323 VGND.n1058 175.546
R2811 VGND.n1729 VGND.n1710 175.546
R2812 VGND.n1727 VGND.n1711 175.546
R2813 VGND.n1716 VGND.n1714 175.546
R2814 VGND.n1068 VGND.n1061 175.546
R2815 VGND.n2007 VGND.n2006 175.546
R2816 VGND.n2014 VGND.n2011 175.546
R2817 VGND.n2020 VGND.n2016 175.546
R2818 VGND.n2027 VGND.n2024 175.546
R2819 VGND.n2025 VGND.n396 175.546
R2820 VGND.n2366 VGND.n1013 175.546
R2821 VGND.n2370 VGND.n2368 175.546
R2822 VGND.n2382 VGND.n1006 175.546
R2823 VGND.n2385 VGND.n2384 175.546
R2824 VGND.n2387 VGND.n1003 175.546
R2825 VGND.n1026 VGND.n1025 175.546
R2826 VGND.n1035 VGND.n1031 175.546
R2827 VGND.n2222 VGND.n2221 175.546
R2828 VGND.n2234 VGND.n2233 175.546
R2829 VGND.n2217 VGND.n2216 175.546
R2830 VGND.n1575 VGND.n997 175.546
R2831 VGND.n2397 VGND.n997 175.546
R2832 VGND.n2397 VGND.n995 175.546
R2833 VGND.n2401 VGND.n995 175.546
R2834 VGND.n2401 VGND.n990 175.546
R2835 VGND.n2412 VGND.n990 175.546
R2836 VGND.n2412 VGND.n988 175.546
R2837 VGND.n2416 VGND.n988 175.546
R2838 VGND.n2416 VGND.n973 175.546
R2839 VGND.n2444 VGND.n973 175.546
R2840 VGND.n2444 VGND.n974 175.546
R2841 VGND.n2711 VGND.n2710 175.546
R2842 VGND.n2708 VGND.n693 175.546
R2843 VGND.n2188 VGND.n2187 175.546
R2844 VGND.n2192 VGND.n984 175.546
R2845 VGND.n2437 VGND.n977 175.546
R2846 VGND.n2990 VGND.n322 175.546
R2847 VGND.n2982 VGND.n2981 175.546
R2848 VGND.n2979 VGND.n332 175.546
R2849 VGND.n2970 VGND.n2969 175.546
R2850 VGND.n2967 VGND.n343 175.546
R2851 VGND.n2849 VGND.n2847 175.546
R2852 VGND.n2808 VGND.n2807 175.546
R2853 VGND.n2810 VGND.n2806 175.546
R2854 VGND.n2789 VGND.n2788 175.546
R2855 VGND.n2791 VGND.n2787 175.546
R2856 VGND.n1803 VGND.n1802 175.546
R2857 VGND.n1808 VGND.n1807 175.546
R2858 VGND.n1817 VGND.n1814 175.546
R2859 VGND.n1822 VGND.n1819 175.546
R2860 VGND.n1824 VGND.n319 175.546
R2861 VGND.n2780 VGND.n2779 175.546
R2862 VGND.n638 VGND.n622 175.546
R2863 VGND.n645 VGND.n640 175.546
R2864 VGND.n643 VGND.n642 175.546
R2865 VGND.n2959 VGND.n352 175.546
R2866 VGND.n2949 VGND.n2948 175.546
R2867 VGND.n2944 VGND.n2943 175.546
R2868 VGND.n2940 VGND.n2939 175.546
R2869 VGND.n604 VGND.n544 175.546
R2870 VGND.n633 VGND.n632 175.546
R2871 VGND.n620 VGND.n616 175.546
R2872 VGND.n611 VGND.n609 175.546
R2873 VGND.n660 VGND.n350 175.546
R2874 VGND.n2545 VGND.n2482 175.546
R2875 VGND.n2541 VGND.n2482 175.546
R2876 VGND.n2541 VGND.n2485 175.546
R2877 VGND.n2490 VGND.n2485 175.546
R2878 VGND.n2530 VGND.n2490 175.546
R2879 VGND.n2530 VGND.n2491 175.546
R2880 VGND.n2526 VGND.n2491 175.546
R2881 VGND.n2526 VGND.n2494 175.546
R2882 VGND.n2519 VGND.n2494 175.546
R2883 VGND.n2519 VGND.n369 175.546
R2884 VGND.n2934 VGND.n369 175.546
R2885 VGND.n2770 VGND.n2769 175.546
R2886 VGND.n2754 VGND.n2753 175.546
R2887 VGND.n2756 VGND.n581 175.546
R2888 VGND.n2480 VGND.n2479 175.546
R2889 VGND.n2549 VGND.n2480 175.546
R2890 VGND.n2706 VGND.n696 175.546
R2891 VGND.n2184 VGND.n697 175.546
R2892 VGND.n2195 VGND.n2194 175.546
R2893 VGND.n2427 VGND.n699 175.546
R2894 VGND.n702 VGND.n699 175.546
R2895 VGND.n2726 VGND.n679 175.546
R2896 VGND.n2141 VGND.n2140 175.546
R2897 VGND.n2136 VGND.n603 175.546
R2898 VGND.n2730 VGND.n595 175.546
R2899 VGND.n674 VGND.n673 175.546
R2900 VGND.n2697 VGND.n706 175.546
R2901 VGND.n2693 VGND.n706 175.546
R2902 VGND.n2693 VGND.n709 175.546
R2903 VGND.n2685 VGND.n709 175.546
R2904 VGND.n2685 VGND.n715 175.546
R2905 VGND.n961 VGND.n715 175.546
R2906 VGND.n2578 VGND.n961 175.546
R2907 VGND.n2578 VGND.n962 175.546
R2908 VGND.n2456 VGND.n962 175.546
R2909 VGND.n2558 VGND.n2456 175.546
R2910 VGND.n2558 VGND.n2457 175.546
R2911 VGND.n582 VGND.n567 175.546
R2912 VGND.n2751 VGND.n572 175.546
R2913 VGND.n2749 VGND.n579 175.546
R2914 VGND.n2471 VGND.n2463 175.546
R2915 VGND.n2461 VGND.n2460 175.546
R2916 VGND.n3027 VGND.n284 175.546
R2917 VGND.n815 VGND.n814 175.546
R2918 VGND.n822 VGND.n817 175.546
R2919 VGND.n820 VGND.n819 175.546
R2920 VGND.n3007 VGND.n312 175.546
R2921 VGND.n1901 VGND.n1899 175.546
R2922 VGND.n1899 VGND.n1654 175.546
R2923 VGND.n1695 VGND.n1654 175.546
R2924 VGND.n1695 VGND.n1658 175.546
R2925 VGND.n1691 VGND.n1658 175.546
R2926 VGND.n1691 VGND.n1660 175.546
R2927 VGND.n1681 VGND.n1660 175.546
R2928 VGND.n1681 VGND.n1666 175.546
R2929 VGND.n1677 VGND.n1666 175.546
R2930 VGND.n1677 VGND.n281 175.546
R2931 VGND.n3030 VGND.n281 175.546
R2932 VGND.n1853 VGND.n1800 175.546
R2933 VGND.n1843 VGND.n1811 175.546
R2934 VGND.n1841 VGND.n1812 175.546
R2935 VGND.n1833 VGND.n1831 175.546
R2936 VGND.n2998 VGND.n317 175.546
R2937 VGND.n1891 VGND.n1753 175.546
R2938 VGND.n1889 VGND.n1754 175.546
R2939 VGND.n1877 VGND.n1776 175.546
R2940 VGND.n1875 VGND.n1777 175.546
R2941 VGND.n1863 VGND.n1860 175.546
R2942 VGND.n2911 VGND.n435 175.546
R2943 VGND.n2909 VGND.n436 175.546
R2944 VGND.n2894 VGND.n2893 175.546
R2945 VGND.n2896 VGND.n2891 175.546
R2946 VGND.n2881 VGND.n2879 175.546
R2947 VGND.n1932 VGND.n1931 175.546
R2948 VGND.n1931 VGND.n1633 175.546
R2949 VGND.n1927 VGND.n1633 175.546
R2950 VGND.n1927 VGND.n1635 175.546
R2951 VGND.n1641 VGND.n1635 175.546
R2952 VGND.n1917 VGND.n1641 175.546
R2953 VGND.n1917 VGND.n1642 175.546
R2954 VGND.n1913 VGND.n1642 175.546
R2955 VGND.n1913 VGND.n1645 175.546
R2956 VGND.n1906 VGND.n1645 175.546
R2957 VGND.n1906 VGND.n1651 175.546
R2958 VGND.n405 VGND.n404 175.546
R2959 VGND.n470 VGND.n407 175.546
R2960 VGND.n473 VGND.n472 175.546
R2961 VGND.n482 VGND.n480 175.546
R2962 VGND.n1797 VGND.n484 175.546
R2963 VGND.n1750 VGND.n1701 175.546
R2964 VGND.n1768 VGND.n1760 175.546
R2965 VGND.n1771 VGND.n1770 175.546
R2966 VGND.n1791 VGND.n1780 175.546
R2967 VGND.n1794 VGND.n1793 175.546
R2968 VGND.n2294 VGND.n2293 175.546
R2969 VGND.n2109 VGND.n2078 175.546
R2970 VGND.n2112 VGND.n2111 175.546
R2971 VGND.n2125 VGND.n2122 175.546
R2972 VGND.n2718 VGND.n684 175.546
R2973 VGND.n2924 VGND.n2923 175.546
R2974 VGND.n2921 VGND.n401 175.546
R2975 VGND.n2866 VGND.n475 175.546
R2976 VGND.n2864 VGND.n476 175.546
R2977 VGND.n2857 VGND.n2856 175.546
R2978 VGND.n2724 VGND.n682 175.546
R2979 VGND.n2150 VGND.n2148 175.546
R2980 VGND.n2146 VGND.n2145 175.546
R2981 VGND.n2738 VGND.n593 175.546
R2982 VGND.n2741 VGND.n2740 175.546
R2983 VGND.n494 VGND.n488 175.546
R2984 VGND.n508 VGND.n499 175.546
R2985 VGND.n511 VGND.n510 175.546
R2986 VGND.n525 VGND.n516 175.546
R2987 VGND.n528 VGND.n527 175.546
R2988 VGND.n589 VGND.n533 175.546
R2989 VGND.n2352 VGND.n1024 175.546
R2990 VGND.n2344 VGND.n2342 175.546
R2991 VGND.n2225 VGND.n2223 175.546
R2992 VGND.n2240 VGND.n2218 175.546
R2993 VGND.n2245 VGND.n2242 175.546
R2994 VGND.n2291 VGND.n2068 175.546
R2995 VGND.n2289 VGND.n2076 175.546
R2996 VGND.n2276 VGND.n2117 175.546
R2997 VGND.n2274 VGND.n2119 175.546
R2998 VGND.n2716 VGND.n687 175.546
R2999 VGND.n1965 VGND.n1964 173.228
R3000 VGND.n1964 VGND.n1963 173.228
R3001 VGND.n1963 VGND.n1601 173.228
R3002 VGND.n1953 VGND.n1601 173.228
R3003 VGND.n1953 VGND.n1952 173.228
R3004 VGND.n1951 VGND.n1609 173.228
R3005 VGND.n1941 VGND.n1609 173.228
R3006 VGND.n1941 VGND.n1940 173.228
R3007 VGND.n1940 VGND.n1939 173.228
R3008 VGND.n1939 VGND.n383 173.228
R3009 VGND.n1930 VGND.n382 173.228
R3010 VGND.n1930 VGND.n1929 173.228
R3011 VGND.n1929 VGND.n1928 173.228
R3012 VGND.n1928 VGND.n1634 173.228
R3013 VGND.n1643 VGND.n1634 173.228
R3014 VGND.n1916 VGND.n1915 173.228
R3015 VGND.n1915 VGND.n1914 173.228
R3016 VGND.n1914 VGND.n1644 173.228
R3017 VGND.n1905 VGND.n1644 173.228
R3018 VGND.n1905 VGND.n1904 173.228
R3019 VGND.n1902 VGND.n1652 173.228
R3020 VGND.n1659 VGND.n1652 173.228
R3021 VGND.n1694 VGND.n1659 173.228
R3022 VGND.n1694 VGND.n1693 173.228
R3023 VGND.n1693 VGND.n1692 173.228
R3024 VGND.n1680 VGND.n1667 173.228
R3025 VGND.n1680 VGND.n1679 173.228
R3026 VGND.n1679 VGND.n1678 173.228
R3027 VGND.n1678 VGND.n280 173.228
R3028 VGND.n3031 VGND.n280 173.228
R3029 VGND.n1204 VGND.n1194 171.863
R3030 VGND.n880 VGND.n879 171.129
R3031 VGND.n913 VGND.n882 171.129
R3032 VGND.n911 VGND.n883 171.129
R3033 VGND.n909 VGND.n885 171.129
R3034 VGND.n907 VGND.n314 171.129
R3035 VGND.n2604 VGND.n810 171.129
R3036 VGND.n2602 VGND.n2601 171.129
R3037 VGND.n859 VGND.n363 171.129
R3038 VGND.n2616 VGND.n797 171.129
R3039 VGND.n868 VGND.n866 171.129
R3040 VGND.n862 VGND.n366 171.129
R3041 VGND.n880 VGND.n869 169.976
R3042 VGND.n914 VGND.n913 169.976
R3043 VGND.n911 VGND.n884 169.976
R3044 VGND.n909 VGND.n886 169.976
R3045 VGND.n907 VGND.n906 169.976
R3046 VGND.n2605 VGND.n2604 169.976
R3047 VGND.n2602 VGND.n804 169.976
R3048 VGND.n935 VGND.n859 169.976
R3049 VGND.n2616 VGND.n2615 169.976
R3050 VGND.n925 VGND.n868 169.976
R3051 VGND.n931 VGND.n862 169.976
R3052 VGND.n879 VGND.n878 168.361
R3053 VGND.n882 VGND.n339 168.361
R3054 VGND.n883 VGND.n328 168.361
R3055 VGND.n885 VGND.n323 168.361
R3056 VGND.n3002 VGND.n314 168.361
R3057 VGND.n810 VGND.n809 168.361
R3058 VGND.n2601 VGND.n835 168.361
R3059 VGND.n797 VGND.n796 168.361
R3060 VGND.n866 VGND.n356 168.361
R3061 VGND.n922 VGND.n869 168.014
R3062 VGND.n914 VGND.n870 168.014
R3063 VGND.n895 VGND.n884 168.014
R3064 VGND.n901 VGND.n886 168.014
R3065 VGND.n906 VGND.n888 168.014
R3066 VGND.n2605 VGND.n805 168.014
R3067 VGND.n2610 VGND.n804 168.014
R3068 VGND.n935 VGND.n934 168.014
R3069 VGND.n2615 VGND.n798 168.014
R3070 VGND.n925 VGND.n924 168.014
R3071 VGND.n932 VGND.n931 168.014
R3072 VGND.t78 VGND.n385 164.887
R3073 VGND.t78 VGND.n386 164.833
R3074 VGND.n2249 VGND.n2248 163.333
R3075 VGND.n2423 VGND.n2422 163.333
R3076 VGND.n2563 VGND.n2562 163.333
R3077 VGND.n1789 VGND.n1788 163.333
R3078 VGND.n3010 VGND.n309 163.333
R3079 VGND.n2886 VGND.n466 163.333
R3080 VGND.n2160 VGND.n2157 163.333
R3081 VGND.n3103 VGND.n199 162.526
R3082 VGND.n1157 VGND.n1091 161.956
R3083 VGND.n1200 VGND.n1199 159.667
R3084 VGND.n1092 VGND.n199 154.468
R3085 VGND.n1157 VGND.n1156 154.315
R3086 VGND.n2510 VGND.n351 153.601
R3087 VGND.n1086 VGND.n1085 152.643
R3088 VGND.n1019 VGND.n1018 152.643
R3089 VGND.n2947 VGND.n2946 152.643
R3090 VGND.n2946 VGND.n2945 152.643
R3091 VGND.n2942 VGND.n2941 152.643
R3092 VGND.n2938 VGND.n2937 152.643
R3093 VGND.n2703 VGND.n2702 152.643
R3094 VGND.n569 VGND.n537 152.643
R3095 VGND.n1164 VGND.n6 152.364
R3096 VGND.n1567 VGND.t91 151.333
R3097 VGND.n1460 VGND.t125 151.333
R3098 VGND.t26 VGND.n3263 151.333
R3099 VGND.n3264 VGND.t26 151.333
R3100 VGND.n2311 VGND.n2310 150
R3101 VGND.n2307 VGND.n2306 150
R3102 VGND.n2303 VGND.n2302 150
R3103 VGND.n2299 VGND.n2298 150
R3104 VGND.n2074 VGND.n2073 150
R3105 VGND.n2286 VGND.n2285 150
R3106 VGND.n2114 VGND.n2113 150
R3107 VGND.n2271 VGND.n2270 150
R3108 VGND.n2348 VGND.n2347 150
R3109 VGND.n2329 VGND.n2328 150
R3110 VGND.n2331 VGND.n1039 150
R3111 VGND.n2236 VGND.n2235 150
R3112 VGND.n2326 VGND.n1055 150
R3113 VGND.n1733 VGND.n1732 150
R3114 VGND.n1724 VGND.n1723 150
R3115 VGND.n1720 VGND.n1719 150
R3116 VGND.n2337 VGND.n2336 150
R3117 VGND.n2339 VGND.n2334 150
R3118 VGND.n2230 VGND.n2228 150
R3119 VGND.n2252 VGND.n2214 150
R3120 VGND.n2254 VGND.n2213 150
R3121 VGND.n2211 VGND.n2210 150
R3122 VGND.n2208 VGND.n2183 150
R3123 VGND.n2425 VGND.n985 150
R3124 VGND.n2394 VGND.n2392 150
R3125 VGND.n2405 VGND.n993 150
R3126 VGND.n2409 VGND.n2407 150
R3127 VGND.n2420 VGND.n986 150
R3128 VGND.n2363 VGND.n2361 150
R3129 VGND.n2375 VGND.n1008 150
R3130 VGND.n2379 VGND.n2377 150
R3131 VGND.n2390 VGND.n1000 150
R3132 VGND.n2201 VGND.n2198 150
R3133 VGND.n2205 VGND.n2203 150
R3134 VGND.n2430 VGND.n981 150
R3135 VGND.n2434 VGND.n2432 150
R3136 VGND.n2260 VGND.n2132 150
R3137 VGND.n2174 VGND.n2172 150
R3138 VGND.n2733 VGND.n601 150
R3139 VGND.n2735 VGND.n600 150
R3140 VGND.n598 VGND.n597 150
R3141 VGND.n2766 VGND.n2765 150
R3142 VGND.n2763 VGND.n577 150
R3143 VGND.n2475 VGND.n2474 150
R3144 VGND.n2690 VGND.n712 150
R3145 VGND.n2688 VGND.n713 150
R3146 VGND.n2573 VGND.n2572 150
R3147 VGND.n2575 VGND.n965 150
R3148 VGND.n2776 VGND.n547 150
R3149 VGND.n635 VGND.n548 150
R3150 VGND.n618 VGND.n617 150
R3151 VGND.n656 VGND.n655 150
R3152 VGND.n573 VGND.n565 150
R3153 VGND.n2760 VGND.n2759 150
R3154 VGND.n2469 VGND.n2468 150
R3155 VGND.n2465 VGND.n2464 150
R3156 VGND.n2538 VGND.n2537 150
R3157 VGND.n2534 VGND.n2533 150
R3158 VGND.n2497 VGND.n2496 150
R3159 VGND.n2523 VGND.n555 150
R3160 VGND.n2516 VGND.n555 150
R3161 VGND.n1756 VGND.n1755 150
R3162 VGND.n1886 VGND.n1885 150
R3163 VGND.n1773 VGND.n1772 150
R3164 VGND.n1872 VGND.n1871 150
R3165 VGND.n425 VGND.n423 150
R3166 VGND.n2918 VGND.n2917 150
R3167 VGND.n477 VGND.n411 150
R3168 VGND.n2861 VGND.n2860 150
R3169 VGND.n2914 VGND.n431 150
R3170 VGND.n445 VGND.n444 150
R3171 VGND.n2900 VGND.n2899 150
R3172 VGND.n462 VGND.n461 150
R3173 VGND.n430 VGND.n422 150
R3174 VGND.n1924 VGND.n422 150
R3175 VGND.n1921 VGND.n1920 150
R3176 VGND.n1647 VGND.n1646 150
R3177 VGND.n1910 VGND.n1909 150
R3178 VGND.n3024 VGND.n3023 150
R3179 VGND.n3021 VGND.n289 150
R3180 VGND.n827 VGND.n826 150
R3181 VGND.n3013 VGND.n3012 150
R3182 VGND.n1848 VGND.n1846 150
R3183 VGND.n1846 VGND.n1805 150
R3184 VGND.n1838 VGND.n1836 150
R3185 VGND.n1828 VGND.n1826 150
R3186 VGND.n1894 VGND.n1699 150
R3187 VGND.n1882 VGND.n1765 150
R3188 VGND.n1880 VGND.n1766 150
R3189 VGND.n1868 VGND.n1785 150
R3190 VGND.n1896 VGND.n1698 150
R3191 VGND.n1686 VGND.n1685 150
R3192 VGND.n1688 VGND.n1684 150
R3193 VGND.n1673 VGND.n1672 150
R3194 VGND.n1674 VGND.n1673 150
R3195 VGND.n2985 VGND.n326 150
R3196 VGND.n2975 VGND.n337 150
R3197 VGND.n2973 VGND.n338 150
R3198 VGND.n2964 VGND.n347 150
R3199 VGND.n628 VGND.n626 150
R3200 VGND.n648 VGND.n614 150
R3201 VGND.n652 VGND.n650 150
R3202 VGND.n2962 VGND.n348 150
R3203 VGND.n2837 VGND.n2836 150
R3204 VGND.n2839 VGND.n2813 150
R3205 VGND.n2796 VGND.n2795 150
R3206 VGND.n2798 VGND.n2794 150
R3207 VGND.n2834 VGND.n2833 150
R3208 VGND.n2833 VGND.n2814 150
R3209 VGND.n2829 VGND.n2827 150
R3210 VGND.n2825 VGND.n2816 150
R3211 VGND.n2821 VGND.n325 150
R3212 VGND.n1623 VGND.n1622 150
R3213 VGND.n2906 VGND.n2905 150
R3214 VGND.n2903 VGND.n443 150
R3215 VGND.n2888 VGND.n465 150
R3216 VGND.n2055 VGND.n2004 150
R3217 VGND.n2047 VGND.n2004 150
R3218 VGND.n2045 VGND.n2013 150
R3219 VGND.n2037 VGND.n2035 150
R3220 VGND.n1972 VGND.n1970 150
R3221 VGND.n1983 VGND.n1076 150
R3222 VGND.n1987 VGND.n1985 150
R3223 VGND.n2001 VGND.n1071 150
R3224 VGND.n1959 VGND.n1605 150
R3225 VGND.n1957 VGND.n1606 150
R3226 VGND.n1947 VGND.n1615 150
R3227 VGND.n1945 VGND.n1616 150
R3228 VGND.n1625 VGND.n1616 150
R3229 VGND.n2844 VGND.n501 150
R3230 VGND.n2842 VGND.n502 150
R3231 VGND.n2803 VGND.n519 150
R3232 VGND.n2801 VGND.n520 150
R3233 VGND.n2264 VGND.n2130 150
R3234 VGND.n2168 VGND.n2155 150
R3235 VGND.n2166 VGND.n2165 150
R3236 VGND.n2163 VGND.n2162 150
R3237 VGND.n2104 VGND.n2103 150
R3238 VGND.n2281 VGND.n2106 150
R3239 VGND.n2279 VGND.n2107 150
R3240 VGND.n2267 VGND.n2129 150
R3241 VGND.n2101 VGND.n2100 150
R3242 VGND.n2100 VGND.n2082 150
R3243 VGND.n2096 VGND.n2094 150
R3244 VGND.n2092 VGND.n2084 150
R3245 VGND.n2088 VGND.n2086 150
R3246 VGND.n136 VGND.n17 146.25
R3247 VGND.n17 VGND.t128 146.25
R3248 VGND.n124 VGND.n18 146.25
R3249 VGND.n18 VGND.t128 146.25
R3250 VGND.n141 VGND.n140 146.25
R3251 VGND.t63 VGND.n141 146.25
R3252 VGND.n130 VGND.n126 146.25
R3253 VGND.t63 VGND.n130 146.25
R3254 VGND.n138 VGND.n118 146.25
R3255 VGND.n118 VGND.t3 146.25
R3256 VGND.n147 VGND.n119 146.25
R3257 VGND.n119 VGND.t3 146.25
R3258 VGND.n24 VGND.n21 146.25
R3259 VGND.t26 VGND.n21 146.25
R3260 VGND.n3260 VGND.n22 146.25
R3261 VGND.t26 VGND.n22 146.25
R3262 VGND.n1596 VGND.n1579 140.875
R3263 VGND.t38 VGND.t60 139.169
R3264 VGND.t60 VGND.t110 139.169
R3265 VGND.t110 VGND.t89 139.169
R3266 VGND.t89 VGND.t115 139.169
R3267 VGND.t55 VGND.t23 139.169
R3268 VGND.t23 VGND.t65 139.169
R3269 VGND.t65 VGND.t40 139.169
R3270 VGND.t40 VGND.t126 139.169
R3271 VGND.n947 VGND.n946 138.204
R3272 VGND.t22 VGND.n384 135.701
R3273 VGND.n3071 VGND.n3070 133.833
R3274 VGND.n1199 VGND.n1198 133.236
R3275 VGND.n3077 VGND.n3076 132.766
R3276 VGND.n2715 VGND.n2714 132.721
R3277 VGND.n1713 VGND.n1712 132.721
R3278 VGND.n2439 VGND.n2438 132.721
R3279 VGND.n536 VGND.n530 132.721
R3280 VGND.n2937 VGND.n2936 132.721
R3281 VGND.n2548 VGND.n2547 132.721
R3282 VGND.n2701 VGND.n2700 132.721
R3283 VGND.n2553 VGND.n586 132.721
R3284 VGND.n2720 VGND.n2719 132.721
R3285 VGND.n3140 VGND.n3139 131.26
R3286 VGND.n1264 VGND.n1172 130.923
R3287 VGND.n104 VGND.n96 127.329
R3288 VGND.n2873 VGND.n387 124.832
R3289 VGND.n876 VGND.n354 124.832
R3290 VGND.n3005 VGND.n313 124.832
R3291 VGND.n1861 VGND.n389 124.832
R3292 VGND.n2931 VGND.n390 124.832
R3293 VGND.n1796 VGND.n388 124.832
R3294 VGND.n3076 VGND.n3075 124.666
R3295 VGND.n3070 VGND.n224 124.543
R3296 VGND.t28 VGND.n782 121.68
R3297 VGND.t68 VGND.n2622 121.68
R3298 VGND.t68 VGND.n769 121.68
R3299 VGND.t13 VGND.n769 121.68
R3300 VGND.t13 VGND.n763 121.68
R3301 VGND.t44 VGND.n763 121.68
R3302 VGND.t30 VGND.n759 121.68
R3303 VGND.t30 VGND.n179 121.68
R3304 VGND.t49 VGND.n179 121.68
R3305 VGND.t49 VGND.n180 121.68
R3306 VGND.t120 VGND.n180 121.68
R3307 VGND.t95 VGND.n161 121.68
R3308 VGND.t94 VGND.n161 121.68
R3309 VGND.t94 VGND.n162 121.68
R3310 VGND.n162 VGND.t96 121.68
R3311 VGND.n3142 VGND.t96 121.68
R3312 VGND.n801 VGND.n800 121.468
R3313 VGND.n3219 VGND.n59 120.77
R3314 VGND.t125 VGND.n1459 117.053
R3315 VGND.n3114 VGND.n3113 117.001
R3316 VGND.t120 VGND.n3114 117.001
R3317 VGND.n3121 VGND.n3120 117.001
R3318 VGND.n3120 VGND.t49 117.001
R3319 VGND.n2656 VGND.n174 117.001
R3320 VGND.t30 VGND.n2656 117.001
R3321 VGND.n2654 VGND.n762 117.001
R3322 VGND.n2654 VGND.t44 117.001
R3323 VGND.n2648 VGND.n2647 117.001
R3324 VGND.t13 VGND.n2648 117.001
R3325 VGND.n2628 VGND.n2627 117.001
R3326 VGND.t68 VGND.n2628 117.001
R3327 VGND.n2633 VGND.n2632 117.001
R3328 VGND.n2632 VGND.t28 117.001
R3329 VGND.n167 VGND.n154 117.001
R3330 VGND.n154 VGND.t96 117.001
R3331 VGND.n3135 VGND.n3134 117.001
R3332 VGND.t94 VGND.n3135 117.001
R3333 VGND.n3110 VGND.n3109 117.001
R3334 VGND.n3109 VGND.t95 117.001
R3335 VGND.n3139 VGND.n155 117.001
R3336 VGND.n155 VGND.t96 117.001
R3337 VGND.n3137 VGND.n3136 117.001
R3338 VGND.n3136 VGND.t94 117.001
R3339 VGND.n3108 VGND.n3107 117.001
R3340 VGND.t95 VGND.n3108 117.001
R3341 VGND.n3116 VGND.n3115 117.001
R3342 VGND.n3115 VGND.t120 117.001
R3343 VGND.n3119 VGND.n3118 117.001
R3344 VGND.t49 VGND.n3119 117.001
R3345 VGND.n2658 VGND.n2657 117.001
R3346 VGND.n2657 VGND.t30 117.001
R3347 VGND.n2653 VGND.n2652 117.001
R3348 VGND.t44 VGND.n2653 117.001
R3349 VGND.n2650 VGND.n2649 117.001
R3350 VGND.n2649 VGND.t13 117.001
R3351 VGND.n2629 VGND.n2621 117.001
R3352 VGND.n2629 VGND.t68 117.001
R3353 VGND.n2631 VGND.n728 117.001
R3354 VGND.t28 VGND.n2631 117.001
R3355 VGND.n1269 VGND.n1161 115.975
R3356 VGND.n106 VGND.n105 115.237
R3357 VGND.n3126 VGND.n156 112.04
R3358 VGND.n1435 VGND.n1434 110.306
R3359 VGND.n1434 VGND.n1433 110.306
R3360 VGND.n1433 VGND.n1432 110.306
R3361 VGND.n1432 VGND.n1431 110.306
R3362 VGND.n1445 VGND.n1392 110.306
R3363 VGND.n1453 VGND.n1392 110.306
R3364 VGND.n1454 VGND.n1453 110.306
R3365 VGND.n1455 VGND.n1454 110.306
R3366 VGND.n2499 VGND.n557 110.023
R3367 VGND.n3034 VGND.n277 109.168
R3368 VGND.n800 VGND.n277 108.433
R3369 VGND.n2505 VGND.n559 106.733
R3370 VGND.n2503 VGND.n560 106.733
R3371 VGND.n2501 VGND.n558 106.733
R3372 VGND.n2501 VGND.n556 106.733
R3373 VGND.n2499 VGND.n556 106.733
R3374 VGND.n2503 VGND.n558 106.733
R3375 VGND.n2505 VGND.n560 106.733
R3376 VGND.t11 VGND.n1311 105.151
R3377 VGND.t11 VGND.n1532 105.151
R3378 VGND.n1532 VGND.t25 105.151
R3379 VGND.n1324 VGND.t25 105.151
R3380 VGND.t32 VGND.n1324 105.151
R3381 VGND.t32 VGND.n1328 105.151
R3382 VGND.t33 VGND.n1328 105.151
R3383 VGND.t33 VGND.n1519 105.151
R3384 VGND.n1519 VGND.t15 105.151
R3385 VGND.n1350 VGND.t15 105.151
R3386 VGND.t5 VGND.n1350 105.151
R3387 VGND.t5 VGND.n1354 105.151
R3388 VGND.t45 VGND.n1354 105.151
R3389 VGND.t45 VGND.n1494 105.151
R3390 VGND.n1494 VGND.t106 105.151
R3391 VGND.n23 VGND.t106 105.151
R3392 VGND.n110 VGND.n109 104.064
R3393 VGND.n1443 VGND.n1435 103.906
R3394 VGND.n1445 VGND.n1444 103.906
R3395 VGND.n1258 VGND.n1257 103.466
R3396 VGND.n1460 VGND.n1311 99.4676
R3397 VGND.n3188 VGND.n3187 97.5005
R3398 VGND.n3187 VGND.n51 97.5005
R3399 VGND.n3157 VGND.n3155 97.5005
R3400 VGND.n3155 VGND.n55 97.5005
R3401 VGND.n3157 VGND.n3156 97.5005
R3402 VGND.n3156 VGND.n90 97.5005
R3403 VGND.n3149 VGND.n3148 97.5005
R3404 VGND.n3148 VGND.n3144 97.5005
R3405 VGND.n3166 VGND.n3165 97.5005
R3406 VGND.n3165 VGND.n51 97.5005
R3407 VGND.n3176 VGND.n3175 97.5005
R3408 VGND.n3175 VGND.n55 97.5005
R3409 VGND.n3176 VGND.n3145 97.5005
R3410 VGND.n3145 VGND.n90 97.5005
R3411 VGND.n3146 VGND.n82 97.5005
R3412 VGND.n3146 VGND.n3144 97.5005
R3413 VGND.n3168 VGND.n3167 97.5005
R3414 VGND.n3167 VGND.n51 97.5005
R3415 VGND.n87 VGND.n86 97.5005
R3416 VGND.n86 VGND.n55 97.5005
R3417 VGND.n88 VGND.n87 97.5005
R3418 VGND.n90 VGND.n88 97.5005
R3419 VGND.n89 VGND.n81 97.5005
R3420 VGND.n3144 VGND.n89 97.5005
R3421 VGND.n116 VGND.n115 97.5005
R3422 VGND.n117 VGND.n116 97.5005
R3423 VGND.n112 VGND.n111 97.5005
R3424 VGND.n111 VGND.n110 97.5005
R3425 VGND.n108 VGND.n97 97.5005
R3426 VGND.n109 VGND.n108 97.5005
R3427 VGND.n104 VGND.n100 97.5005
R3428 VGND.n100 VGND.n99 97.5005
R3429 VGND.n66 VGND.n49 97.5005
R3430 VGND.n51 VGND.n49 97.5005
R3431 VGND.n62 VGND.n50 97.5005
R3432 VGND.n55 VGND.n50 97.5005
R3433 VGND.n3213 VGND.n62 97.5005
R3434 VGND.n3213 VGND.n90 97.5005
R3435 VGND.n3220 VGND.n3219 97.5005
R3436 VGND.n3220 VGND.n3144 97.5005
R3437 VGND.n3267 VGND.n3266 97.5005
R3438 VGND.n3268 VGND.n3267 97.5005
R3439 VGND.n133 VGND.n132 97.5005
R3440 VGND.n132 VGND.n131 97.5005
R3441 VGND.n134 VGND.n133 97.5005
R3442 VGND.n134 VGND.n129 97.5005
R3443 VGND.n145 VGND.n128 97.5005
R3444 VGND.n142 VGND.n128 97.5005
R3445 VGND.n145 VGND.n144 97.5005
R3446 VGND.n144 VGND.n143 97.5005
R3447 VGND.n149 VGND.n148 97.5005
R3448 VGND.n150 VGND.n149 97.5005
R3449 VGND.n3262 VGND.n3261 97.5005
R3450 VGND.n3263 VGND.n3262 97.5005
R3451 VGND.n3266 VGND.n3265 97.5005
R3452 VGND.n3265 VGND.n3264 97.5005
R3453 VGND.n1431 VGND.n1382 97.5005
R3454 VGND.t76 VGND.n1382 97.5005
R3455 VGND.n1433 VGND.n1395 97.5005
R3456 VGND.t51 VGND.n1395 97.5005
R3457 VGND.n1435 VGND.n1402 97.5005
R3458 VGND.t98 VGND.n1402 97.5005
R3459 VGND.n1467 VGND.n1466 97.5005
R3460 VGND.n1466 VGND.t76 97.5005
R3461 VGND.n1416 VGND.n1396 97.5005
R3462 VGND.t51 VGND.n1396 97.5005
R3463 VGND.n1406 VGND.n1403 97.5005
R3464 VGND.t98 VGND.n1403 97.5005
R3465 VGND.n1465 VGND.n1464 97.5005
R3466 VGND.t76 VGND.n1465 97.5005
R3467 VGND.n1451 VGND.n1450 97.5005
R3468 VGND.t51 VGND.n1451 97.5005
R3469 VGND.n1448 VGND.n1447 97.5005
R3470 VGND.n1447 VGND.t98 97.5005
R3471 VGND.n1455 VGND.n1383 97.5005
R3472 VGND.t76 VGND.n1383 97.5005
R3473 VGND.n1453 VGND.n1452 97.5005
R3474 VGND.n1452 VGND.t51 97.5005
R3475 VGND.n1446 VGND.n1445 97.5005
R3476 VGND.t98 VGND.n1446 97.5005
R3477 VGND.t52 VGND.n380 96.247
R3478 VGND.n1498 VGND.n1497 94.3594
R3479 VGND.n1189 VGND.n1165 94.255
R3480 VGND.t120 VGND.n188 93.6388
R3481 VGND.n3272 VGND.n13 93.538
R3482 VGND.n2728 VGND.t78 92.209
R3483 VGND.n399 VGND.t78 92.209
R3484 VGND.n1952 VGND.t78 90.4642
R3485 VGND.t78 VGND.n1643 90.4642
R3486 VGND.n1692 VGND.t78 90.4642
R3487 VGND.n3268 VGND.t128 90.0553
R3488 VGND.n131 VGND.t128 90.0553
R3489 VGND.t63 VGND.n129 90.0553
R3490 VGND.n142 VGND.t63 90.0553
R3491 VGND.n143 VGND.t3 90.0553
R3492 VGND.n1431 VGND.n1390 89.224
R3493 VGND.n1456 VGND.n1455 89.224
R3494 VGND.n25 VGND.t27 88.4435
R3495 VGND.n120 VGND.t64 88.4111
R3496 VGND.n3245 VGND.t119 88.0285
R3497 VGND.n3160 VGND.t117 88.0261
R3498 VGND.n3151 VGND.t67 88.0261
R3499 VGND.n3180 VGND.t92 87.9901
R3500 VGND.n3174 VGND.t73 87.9901
R3501 VGND.n3194 VGND.t75 87.9804
R3502 VGND.n3195 VGND.t36 87.9804
R3503 VGND.n31 VGND.t43 87.9324
R3504 VGND.n3232 VGND.t113 87.9252
R3505 VGND.n64 VGND.t47 87.9252
R3506 VGND.n2442 VGND.n2441 87.7399
R3507 VGND.n2556 VGND.n2555 87.7399
R3508 VGND.n25 VGND.t129 87.5033
R3509 VGND.n120 VGND.t4 87.4792
R3510 VGND.n151 VGND.t3 87.0957
R3511 VGND.n3236 VGND.n59 84.9783
R3512 VGND.n1497 VGND.n12 83.9475
R3513 VGND.n3237 VGND.n3236 83.7931
R3514 VGND.n2696 VGND.n707 83.3964
R3515 VGND.n2544 VGND.n2481 83.3964
R3516 VGND.t44 VGND.t6 83.1233
R3517 VGND.t78 VGND.n1951 82.7652
R3518 VGND.n1916 VGND.t78 82.7652
R3519 VGND.n1667 VGND.t78 82.7652
R3520 VGND.n3273 VGND.n3272 82.7361
R3521 VGND.n1184 VGND.n1176 80.2978
R3522 VGND.t11 VGND.n1315 79.8338
R3523 VGND.t11 VGND.n1312 79.8338
R3524 VGND.t25 VGND.n1312 79.8338
R3525 VGND.n1327 VGND.t25 79.8338
R3526 VGND.t32 VGND.n1327 79.8338
R3527 VGND.t32 VGND.n1325 79.8338
R3528 VGND.t33 VGND.n1325 79.8338
R3529 VGND.t33 VGND.n1339 79.8338
R3530 VGND.t15 VGND.n1339 79.8338
R3531 VGND.n1353 VGND.t15 79.8338
R3532 VGND.t5 VGND.n1353 79.8338
R3533 VGND.t5 VGND.n1351 79.8338
R3534 VGND.t45 VGND.n1351 79.8338
R3535 VGND.t45 VGND.n1367 79.8338
R3536 VGND.n1367 VGND.t106 79.8338
R3537 VGND.n3270 VGND.t106 79.8338
R3538 VGND.n1587 VGND.n1586 78.7861
R3539 VGND.n2582 VGND.n719 78.6088
R3540 VGND.n1576 VGND.n996 78.1841
R3541 VGND.n2398 VGND.n996 78.1841
R3542 VGND.n2399 VGND.n2398 78.1841
R3543 VGND.n2400 VGND.n2399 78.1841
R3544 VGND.n2400 VGND.n989 78.1841
R3545 VGND.n2413 VGND.n989 78.1841
R3546 VGND.n2414 VGND.n2413 78.1841
R3547 VGND.n2415 VGND.n2414 78.1841
R3548 VGND.n2415 VGND.n975 78.1841
R3549 VGND.n2443 VGND.n975 78.1841
R3550 VGND.n2443 VGND.n2442 78.1841
R3551 VGND.n2696 VGND.n2695 78.1841
R3552 VGND.n2695 VGND.n2694 78.1841
R3553 VGND.n2694 VGND.n708 78.1841
R3554 VGND.n2684 VGND.n708 78.1841
R3555 VGND.n2684 VGND.n2683 78.1841
R3556 VGND.n2579 VGND.n959 78.1841
R3557 VGND.n2458 VGND.n959 78.1841
R3558 VGND.n2557 VGND.n2458 78.1841
R3559 VGND.n2557 VGND.n2556 78.1841
R3560 VGND.n2544 VGND.n2543 78.1841
R3561 VGND.n2543 VGND.n2542 78.1841
R3562 VGND.n2542 VGND.n2484 78.1841
R3563 VGND.n2492 VGND.n2484 78.1841
R3564 VGND.n2529 VGND.n2492 78.1841
R3565 VGND.n2529 VGND.n2528 78.1841
R3566 VGND.n2528 VGND.n2527 78.1841
R3567 VGND.n2527 VGND.n2493 78.1841
R3568 VGND.n2518 VGND.n2493 78.1841
R3569 VGND.n2518 VGND.n371 78.1841
R3570 VGND.n2933 VGND.n371 78.1841
R3571 VGND.n3202 VGND.n3201 76.8427
R3572 VGND.n1087 VGND.n1086 76.3222
R3573 VGND.n1977 VGND.n1976 76.3222
R3574 VGND.n1980 VGND.n1979 76.3222
R3575 VGND.n1992 VGND.n1991 76.3222
R3576 VGND.n1998 VGND.n1997 76.3222
R3577 VGND.n1631 VGND.n1630 76.3222
R3578 VGND.n439 VGND.n438 76.3222
R3579 VGND.n453 VGND.n452 76.3222
R3580 VGND.n456 VGND.n455 76.3222
R3581 VGND.n2877 VGND.n2876 76.3222
R3582 VGND.n2874 VGND.n2873 76.3222
R3583 VGND.n2062 VGND.n2061 76.3222
R3584 VGND.n2051 VGND.n1067 76.3222
R3585 VGND.n2050 VGND.n2009 76.3222
R3586 VGND.n2042 VGND.n2041 76.3222
R3587 VGND.n2031 VGND.n2018 76.3222
R3588 VGND.n2030 VGND.n2029 76.3222
R3589 VGND.n2319 VGND.n2318 76.3222
R3590 VGND.n2322 VGND.n2321 76.3222
R3591 VGND.n1709 VGND.n1058 76.3222
R3592 VGND.n1729 VGND.n1728 76.3222
R3593 VGND.n1715 VGND.n1711 76.3222
R3594 VGND.n1714 VGND.n1713 76.3222
R3595 VGND.n2006 VGND.n2005 76.3222
R3596 VGND.n2011 VGND.n2010 76.3222
R3597 VGND.n2016 VGND.n2015 76.3222
R3598 VGND.n2024 VGND.n2023 76.3222
R3599 VGND.n2026 VGND.n2025 76.3222
R3600 VGND.n1020 VGND.n1019 76.3222
R3601 VGND.n2367 VGND.n2366 76.3222
R3602 VGND.n2370 VGND.n2369 76.3222
R3603 VGND.n2383 VGND.n2382 76.3222
R3604 VGND.n2386 VGND.n2385 76.3222
R3605 VGND.n1025 VGND.n672 76.3222
R3606 VGND.n1031 VGND.n671 76.3222
R3607 VGND.n2221 VGND.n670 76.3222
R3608 VGND.n2233 VGND.n669 76.3222
R3609 VGND.n2216 VGND.n668 76.3222
R3610 VGND.n690 VGND.n667 76.3222
R3611 VGND.n2712 VGND.n2711 76.3222
R3612 VGND.n2709 VGND.n2708 76.3222
R3613 VGND.n2187 VGND.n2186 76.3222
R3614 VGND.n2192 VGND.n2191 76.3222
R3615 VGND.n983 VGND.n977 76.3222
R3616 VGND.n2991 VGND.n2990 76.3222
R3617 VGND.n2982 VGND.n329 76.3222
R3618 VGND.n2980 VGND.n2979 76.3222
R3619 VGND.n2970 VGND.n340 76.3222
R3620 VGND.n2968 VGND.n2967 76.3222
R3621 VGND.n876 VGND.n875 76.3222
R3622 VGND.n2848 VGND.n491 76.3222
R3623 VGND.n2847 VGND.n496 76.3222
R3624 VGND.n2809 VGND.n2808 76.3222
R3625 VGND.n2806 VGND.n513 76.3222
R3626 VGND.n2790 VGND.n2789 76.3222
R3627 VGND.n2787 VGND.n530 76.3222
R3628 VGND.n1802 VGND.n1801 76.3222
R3629 VGND.n1807 VGND.n1806 76.3222
R3630 VGND.n1814 VGND.n1813 76.3222
R3631 VGND.n1819 VGND.n1818 76.3222
R3632 VGND.n1824 VGND.n1823 76.3222
R3633 VGND.n2993 VGND.n321 76.3222
R3634 VGND.n2782 VGND.n2781 76.3222
R3635 VGND.n2779 VGND.n542 76.3222
R3636 VGND.n639 VGND.n638 76.3222
R3637 VGND.n645 VGND.n644 76.3222
R3638 VGND.n642 VGND.n641 76.3222
R3639 VGND.n2958 VGND.n2957 76.3222
R3640 VGND.n2949 VGND.n368 76.3222
R3641 VGND.n2945 VGND.n2944 76.3222
R3642 VGND.n2941 VGND.n2940 76.3222
R3643 VGND.n605 VGND.n604 76.3222
R3644 VGND.n632 VGND.n606 76.3222
R3645 VGND.n620 VGND.n607 76.3222
R3646 VGND.n611 VGND.n608 76.3222
R3647 VGND.n661 VGND.n660 76.3222
R3648 VGND.n666 VGND.n665 76.3222
R3649 VGND.n538 VGND.n537 76.3222
R3650 VGND.n2770 VGND.n569 76.3222
R3651 VGND.n2769 VGND.n570 76.3222
R3652 VGND.n2755 VGND.n2754 76.3222
R3653 VGND.n2478 VGND.n581 76.3222
R3654 VGND.n2702 VGND.n698 76.3222
R3655 VGND.n2703 VGND.n696 76.3222
R3656 VGND.n2706 VGND.n2705 76.3222
R3657 VGND.n2184 VGND.n701 76.3222
R3658 VGND.n2194 VGND.n700 76.3222
R3659 VGND.n2727 VGND.n2726 76.3222
R3660 VGND.n2141 VGND.n677 76.3222
R3661 VGND.n2136 VGND.n676 76.3222
R3662 VGND.n2730 VGND.n2729 76.3222
R3663 VGND.n675 VGND.n674 76.3222
R3664 VGND.n2745 VGND.n587 76.3222
R3665 VGND.n2746 VGND.n582 76.3222
R3666 VGND.n583 VGND.n572 76.3222
R3667 VGND.n2750 VGND.n2749 76.3222
R3668 VGND.n2471 VGND.n584 76.3222
R3669 VGND.n2460 VGND.n585 76.3222
R3670 VGND.n3028 VGND.n3027 76.3222
R3671 VGND.n814 VGND.n813 76.3222
R3672 VGND.n817 VGND.n816 76.3222
R3673 VGND.n821 VGND.n820 76.3222
R3674 VGND.n818 VGND.n312 76.3222
R3675 VGND.n3006 VGND.n3005 76.3222
R3676 VGND.n1855 VGND.n1854 76.3222
R3677 VGND.n1810 VGND.n1800 76.3222
R3678 VGND.n1843 VGND.n1842 76.3222
R3679 VGND.n1832 VGND.n1812 76.3222
R3680 VGND.n1831 VGND.n1821 76.3222
R3681 VGND.n2999 VGND.n2998 76.3222
R3682 VGND.n1752 VGND.n1653 76.3222
R3683 VGND.n1891 VGND.n1890 76.3222
R3684 VGND.n1775 VGND.n1754 76.3222
R3685 VGND.n1877 VGND.n1876 76.3222
R3686 VGND.n1859 VGND.n1777 76.3222
R3687 VGND.n1863 VGND.n1862 76.3222
R3688 VGND.n1934 VGND.n1933 76.3222
R3689 VGND.n2911 VGND.n2910 76.3222
R3690 VGND.n2892 VGND.n436 76.3222
R3691 VGND.n2895 VGND.n2894 76.3222
R3692 VGND.n2891 VGND.n458 76.3222
R3693 VGND.n2881 VGND.n2880 76.3222
R3694 VGND.n404 VGND.n403 76.3222
R3695 VGND.n406 VGND.n405 76.3222
R3696 VGND.n471 VGND.n470 76.3222
R3697 VGND.n479 VGND.n473 76.3222
R3698 VGND.n483 VGND.n482 76.3222
R3699 VGND.n1798 VGND.n1797 76.3222
R3700 VGND.n1749 VGND.n1748 76.3222
R3701 VGND.n1759 VGND.n1701 76.3222
R3702 VGND.n1769 VGND.n1768 76.3222
R3703 VGND.n1779 VGND.n1771 76.3222
R3704 VGND.n1792 VGND.n1791 76.3222
R3705 VGND.n1795 VGND.n1794 76.3222
R3706 VGND.n1796 VGND.n1795 76.3222
R3707 VGND.n1793 VGND.n1792 76.3222
R3708 VGND.n1780 VGND.n1779 76.3222
R3709 VGND.n1770 VGND.n1769 76.3222
R3710 VGND.n1760 VGND.n1759 76.3222
R3711 VGND.n1750 VGND.n1749 76.3222
R3712 VGND.n1753 VGND.n1752 76.3222
R3713 VGND.n1890 VGND.n1889 76.3222
R3714 VGND.n1776 VGND.n1775 76.3222
R3715 VGND.n1876 VGND.n1875 76.3222
R3716 VGND.n1860 VGND.n1859 76.3222
R3717 VGND.n1862 VGND.n1861 76.3222
R3718 VGND.n321 VGND.n319 76.3222
R3719 VGND.n1823 VGND.n1822 76.3222
R3720 VGND.n1818 VGND.n1817 76.3222
R3721 VGND.n1813 VGND.n1808 76.3222
R3722 VGND.n1806 VGND.n1803 76.3222
R3723 VGND.n1801 VGND.n490 76.3222
R3724 VGND.n407 VGND.n406 76.3222
R3725 VGND.n472 VGND.n471 76.3222
R3726 VGND.n480 VGND.n479 76.3222
R3727 VGND.n484 VGND.n483 76.3222
R3728 VGND.n1799 VGND.n1798 76.3222
R3729 VGND.n1854 VGND.n1853 76.3222
R3730 VGND.n1811 VGND.n1810 76.3222
R3731 VGND.n1842 VGND.n1841 76.3222
R3732 VGND.n1833 VGND.n1832 76.3222
R3733 VGND.n1821 VGND.n317 76.3222
R3734 VGND.n3000 VGND.n2999 76.3222
R3735 VGND.n2939 VGND.n2938 76.3222
R3736 VGND.n2943 VGND.n2942 76.3222
R3737 VGND.n2948 VGND.n2947 76.3222
R3738 VGND.n662 VGND.n368 76.3222
R3739 VGND.n875 VGND.n343 76.3222
R3740 VGND.n2969 VGND.n2968 76.3222
R3741 VGND.n340 VGND.n332 76.3222
R3742 VGND.n2981 VGND.n2980 76.3222
R3743 VGND.n329 VGND.n322 76.3222
R3744 VGND.n2992 VGND.n2991 76.3222
R3745 VGND.n3007 VGND.n3006 76.3222
R3746 VGND.n819 VGND.n818 76.3222
R3747 VGND.n822 VGND.n821 76.3222
R3748 VGND.n816 VGND.n815 76.3222
R3749 VGND.n813 VGND.n284 76.3222
R3750 VGND.n3029 VGND.n3028 76.3222
R3751 VGND.n2438 VGND.n2437 76.3222
R3752 VGND.n984 VGND.n983 76.3222
R3753 VGND.n2191 VGND.n2188 76.3222
R3754 VGND.n2186 VGND.n693 76.3222
R3755 VGND.n2710 VGND.n2709 76.3222
R3756 VGND.n2705 VGND.n697 76.3222
R3757 VGND.n2195 VGND.n701 76.3222
R3758 VGND.n2427 VGND.n700 76.3222
R3759 VGND.n2701 VGND.n702 76.3222
R3760 VGND.n2027 VGND.n2026 76.3222
R3761 VGND.n2023 VGND.n2020 76.3222
R3762 VGND.n2015 VGND.n2014 76.3222
R3763 VGND.n2010 VGND.n2007 76.3222
R3764 VGND.n2005 VGND.n1068 76.3222
R3765 VGND.n2061 VGND.n2060 76.3222
R3766 VGND.n2052 VGND.n2051 76.3222
R3767 VGND.n2017 VGND.n2009 76.3222
R3768 VGND.n2041 VGND.n2040 76.3222
R3769 VGND.n2032 VGND.n2031 76.3222
R3770 VGND.n2294 VGND.n2070 76.3222
R3771 VGND.n2293 VGND.n2071 76.3222
R3772 VGND.n2110 VGND.n2109 76.3222
R3773 VGND.n2121 VGND.n2112 76.3222
R3774 VGND.n2125 VGND.n2124 76.3222
R3775 VGND.n2719 VGND.n2718 76.3222
R3776 VGND.n2078 VGND.n2071 76.3222
R3777 VGND.n2111 VGND.n2110 76.3222
R3778 VGND.n2122 VGND.n2121 76.3222
R3779 VGND.n2124 VGND.n684 76.3222
R3780 VGND.n2925 VGND.n2924 76.3222
R3781 VGND.n2922 VGND.n2921 76.3222
R3782 VGND.n475 VGND.n474 76.3222
R3783 VGND.n2865 VGND.n2864 76.3222
R3784 VGND.n2857 VGND.n486 76.3222
R3785 VGND.n2855 VGND.n2854 76.3222
R3786 VGND.n2856 VGND.n2855 76.3222
R3787 VGND.n486 VGND.n476 76.3222
R3788 VGND.n2866 VGND.n2865 76.3222
R3789 VGND.n474 VGND.n401 76.3222
R3790 VGND.n2923 VGND.n2922 76.3222
R3791 VGND.n2723 VGND.n2722 76.3222
R3792 VGND.n2149 VGND.n682 76.3222
R3793 VGND.n2148 VGND.n2147 76.3222
R3794 VGND.n2145 VGND.n2142 76.3222
R3795 VGND.n2739 VGND.n2738 76.3222
R3796 VGND.n2742 VGND.n2741 76.3222
R3797 VGND.n499 VGND.n498 76.3222
R3798 VGND.n510 VGND.n509 76.3222
R3799 VGND.n516 VGND.n515 76.3222
R3800 VGND.n527 VGND.n526 76.3222
R3801 VGND.n533 VGND.n532 76.3222
R3802 VGND.n532 VGND.n528 76.3222
R3803 VGND.n526 VGND.n525 76.3222
R3804 VGND.n515 VGND.n511 76.3222
R3805 VGND.n509 VGND.n508 76.3222
R3806 VGND.n498 VGND.n494 76.3222
R3807 VGND.n2849 VGND.n2848 76.3222
R3808 VGND.n2807 VGND.n496 76.3222
R3809 VGND.n2810 VGND.n2809 76.3222
R3810 VGND.n2788 VGND.n513 76.3222
R3811 VGND.n2791 VGND.n2790 76.3222
R3812 VGND.n2461 VGND.n586 76.3222
R3813 VGND.n2463 VGND.n585 76.3222
R3814 VGND.n584 VGND.n579 76.3222
R3815 VGND.n2751 VGND.n2750 76.3222
R3816 VGND.n583 VGND.n567 76.3222
R3817 VGND.n2753 VGND.n570 76.3222
R3818 VGND.n2756 VGND.n2755 76.3222
R3819 VGND.n2479 VGND.n2478 76.3222
R3820 VGND.n2549 VGND.n2548 76.3222
R3821 VGND.n2217 VGND.n667 76.3222
R3822 VGND.n2234 VGND.n668 76.3222
R3823 VGND.n2222 VGND.n669 76.3222
R3824 VGND.n1035 VGND.n670 76.3222
R3825 VGND.n1026 VGND.n671 76.3222
R3826 VGND.n1021 VGND.n672 76.3222
R3827 VGND.n2712 VGND.n691 76.3222
R3828 VGND.n673 VGND.n587 76.3222
R3829 VGND.n675 VGND.n595 76.3222
R3830 VGND.n2729 VGND.n603 76.3222
R3831 VGND.n2140 VGND.n676 76.3222
R3832 VGND.n679 VGND.n677 76.3222
R3833 VGND.n2727 VGND.n678 76.3222
R3834 VGND.n2747 VGND.n2746 76.3222
R3835 VGND.n666 VGND.n350 76.3222
R3836 VGND.n661 VGND.n609 76.3222
R3837 VGND.n616 VGND.n608 76.3222
R3838 VGND.n633 VGND.n607 76.3222
R3839 VGND.n606 VGND.n544 76.3222
R3840 VGND.n605 VGND.n539 76.3222
R3841 VGND.n2724 VGND.n2723 76.3222
R3842 VGND.n2150 VGND.n2149 76.3222
R3843 VGND.n2147 VGND.n2146 76.3222
R3844 VGND.n2142 VGND.n593 76.3222
R3845 VGND.n2740 VGND.n2739 76.3222
R3846 VGND.n2743 VGND.n2742 76.3222
R3847 VGND.n2781 VGND.n2780 76.3222
R3848 VGND.n622 VGND.n542 76.3222
R3849 VGND.n640 VGND.n639 76.3222
R3850 VGND.n644 VGND.n643 76.3222
R3851 VGND.n641 VGND.n352 76.3222
R3852 VGND.n2959 VGND.n2958 76.3222
R3853 VGND.n2354 VGND.n2353 76.3222
R3854 VGND.n2343 VGND.n1024 76.3222
R3855 VGND.n2342 VGND.n1033 76.3222
R3856 VGND.n2225 VGND.n2224 76.3222
R3857 VGND.n2241 VGND.n2240 76.3222
R3858 VGND.n2245 VGND.n2244 76.3222
R3859 VGND.n2353 VGND.n2352 76.3222
R3860 VGND.n2344 VGND.n2343 76.3222
R3861 VGND.n2223 VGND.n1033 76.3222
R3862 VGND.n2224 VGND.n2218 76.3222
R3863 VGND.n2242 VGND.n2241 76.3222
R3864 VGND.n2244 VGND.n2243 76.3222
R3865 VGND.n2068 VGND.n2067 76.3222
R3866 VGND.n2290 VGND.n2289 76.3222
R3867 VGND.n2117 VGND.n2116 76.3222
R3868 VGND.n2275 VGND.n2274 76.3222
R3869 VGND.n2118 VGND.n687 76.3222
R3870 VGND.n2716 VGND.n2715 76.3222
R3871 VGND.n2119 VGND.n2118 76.3222
R3872 VGND.n2276 VGND.n2275 76.3222
R3873 VGND.n2116 VGND.n2076 76.3222
R3874 VGND.n2291 VGND.n2290 76.3222
R3875 VGND.n2067 VGND.n2066 76.3222
R3876 VGND.n2070 VGND.n398 76.3222
R3877 VGND.n2926 VGND.n2925 76.3222
R3878 VGND.n2029 VGND.n393 76.3222
R3879 VGND.n403 VGND.n391 76.3222
R3880 VGND.n2875 VGND.n2874 76.3222
R3881 VGND.n2876 VGND.n460 76.3222
R3882 VGND.n455 VGND.n454 76.3222
R3883 VGND.n452 VGND.n451 76.3222
R3884 VGND.n438 VGND.n433 76.3222
R3885 VGND.n1630 VGND.n1629 76.3222
R3886 VGND.n1933 VGND.n435 76.3222
R3887 VGND.n2910 VGND.n2909 76.3222
R3888 VGND.n2893 VGND.n2892 76.3222
R3889 VGND.n2896 VGND.n2895 76.3222
R3890 VGND.n2879 VGND.n458 76.3222
R3891 VGND.n2880 VGND.n390 76.3222
R3892 VGND.n1018 VGND.n1013 76.3222
R3893 VGND.n2368 VGND.n2367 76.3222
R3894 VGND.n2369 VGND.n1006 76.3222
R3895 VGND.n2384 VGND.n2383 76.3222
R3896 VGND.n2387 VGND.n2386 76.3222
R3897 VGND.n2320 VGND.n2319 76.3222
R3898 VGND.n2323 VGND.n2322 76.3222
R3899 VGND.n1710 VGND.n1709 76.3222
R3900 VGND.n1728 VGND.n1727 76.3222
R3901 VGND.n1716 VGND.n1715 76.3222
R3902 VGND.n1085 VGND.n1080 76.3222
R3903 VGND.n1978 VGND.n1977 76.3222
R3904 VGND.n1979 VGND.n1073 76.3222
R3905 VGND.n1993 VGND.n1992 76.3222
R3906 VGND.n1997 VGND.n1996 76.3222
R3907 VGND.n2915 VGND.n2914 76.062
R3908 VGND.n1895 VGND.n1894 76.062
R3909 VGND.n1896 VGND.n1895 76.062
R3910 VGND.n2915 VGND.n430 76.062
R3911 VGND.n2836 VGND.n2835 76.062
R3912 VGND.n2835 VGND.n2834 76.062
R3913 VGND.n1970 VGND.n1082 76.062
R3914 VGND.n1605 VGND.n1082 76.062
R3915 VGND.n2103 VGND.n2102 76.062
R3916 VGND.n2102 VGND.n2101 76.062
R3917 VGND.n2298 VGND.n1044 74.5978
R3918 VGND.n2253 VGND.n2252 74.5978
R3919 VGND.n600 VGND.n599 74.5978
R3920 VGND.n1755 VGND.n412 74.5978
R3921 VGND.n3024 VGND.n287 74.5978
R3922 VGND.n1674 VGND.n287 74.5978
R3923 VGND.n1909 VGND.n412 74.5978
R3924 VGND.n2254 VGND.n2253 74.5978
R3925 VGND.n1624 VGND.n1623 74.5978
R3926 VGND.n1625 VGND.n1624 74.5978
R3927 VGND.n2086 VGND.n2085 74.5978
R3928 VGND.n2073 VGND.n1044 74.5978
R3929 VGND.n2085 VGND.n501 74.5978
R3930 VGND.n599 VGND.n598 74.5978
R3931 VGND.n1459 VGND.n1315 73.3608
R3932 VGND.t28 VGND.n2619 72.6078
R3933 VGND.n2513 VGND.n2512 71.7719
R3934 VGND.n2512 VGND.n2511 70.4005
R3935 VGND.n2511 VGND.n2510 69.9434
R3936 VGND.n1266 VGND.t115 69.5849
R3937 VGND.n2348 VGND.n1028 69.3109
R3938 VGND.n2392 VGND.n2391 69.3109
R3939 VGND.n2434 VGND.n2433 69.3109
R3940 VGND.n2464 VGND.n561 69.3109
R3941 VGND.n2537 VGND.n561 69.3109
R3942 VGND.n2391 VGND.n2390 69.3109
R3943 VGND.n2433 VGND.n712 69.3109
R3944 VGND.n1719 VGND.n1028 69.3109
R3945 VGND.n707 VGND.t78 68.6283
R3946 VGND.n2481 VGND.t78 68.6283
R3947 VGND.n1588 VGND.n1580 67.7944
R3948 VGND.n2441 VGND.t78 67.7596
R3949 VGND.n2555 VGND.t78 67.7596
R3950 VGND.n3035 VGND.n276 66.8968
R3951 VGND.n3259 VGND.n24 66.8643
R3952 VGND.n1457 VGND.n1456 65.8695
R3953 VGND.n2504 VGND.n2503 65.8183
R3954 VGND.t79 VGND.n560 65.8183
R3955 VGND.n2506 VGND.n2505 65.8183
R3956 VGND.t79 VGND.n559 65.8183
R3957 VGND.n2502 VGND.n2501 65.8183
R3958 VGND.t79 VGND.n558 65.8183
R3959 VGND.n2500 VGND.n2499 65.8183
R3960 VGND.t79 VGND.n556 65.8183
R3961 VGND.t84 VGND.n417 65.8183
R3962 VGND.t84 VGND.n419 65.8183
R3963 VGND.n2916 VGND.t84 65.8183
R3964 VGND.t84 VGND.n409 65.8183
R3965 VGND.n1664 VGND.t82 65.8183
R3966 VGND.n1687 VGND.t82 65.8183
R3967 VGND.n1656 VGND.t82 65.8183
R3968 VGND.t84 VGND.n418 65.8183
R3969 VGND.t84 VGND.n420 65.8183
R3970 VGND.t84 VGND.n421 65.8183
R3971 VGND.t84 VGND.n416 65.8183
R3972 VGND.t84 VGND.n415 65.8183
R3973 VGND.t84 VGND.n414 65.8183
R3974 VGND.t84 VGND.n413 65.8183
R3975 VGND.n1764 VGND.t82 65.8183
R3976 VGND.n1881 VGND.t82 65.8183
R3977 VGND.n1784 VGND.t82 65.8183
R3978 VGND.n1867 VGND.t82 65.8183
R3979 VGND.n1827 VGND.t82 65.8183
R3980 VGND.n1815 VGND.t82 65.8183
R3981 VGND.n1837 VGND.t82 65.8183
R3982 VGND.n1847 VGND.t82 65.8183
R3983 VGND.n3011 VGND.t82 65.8183
R3984 VGND.n307 VGND.t82 65.8183
R3985 VGND.n824 VGND.t82 65.8183
R3986 VGND.n3022 VGND.t82 65.8183
R3987 VGND.n346 VGND.t85 65.8183
R3988 VGND.n2974 VGND.t85 65.8183
R3989 VGND.n335 VGND.t85 65.8183
R3990 VGND.n2986 VGND.t85 65.8183
R3991 VGND.n2820 VGND.t85 65.8183
R3992 VGND.n2826 VGND.t85 65.8183
R3993 VGND.n2828 VGND.t85 65.8183
R3994 VGND.n2561 VGND.t80 65.8183
R3995 VGND.n2574 VGND.t80 65.8183
R3996 VGND.n2571 VGND.t80 65.8183
R3997 VGND.t79 VGND.n553 65.8183
R3998 VGND.t79 VGND.n551 65.8183
R3999 VGND.t79 VGND.n549 65.8183
R4000 VGND.n2360 VGND.t86 65.8183
R4001 VGND.n2362 VGND.t86 65.8183
R4002 VGND.n2376 VGND.t86 65.8183
R4003 VGND.n2378 VGND.t86 65.8183
R4004 VGND.n2421 VGND.t86 65.8183
R4005 VGND.n2408 VGND.t86 65.8183
R4006 VGND.n2406 VGND.t86 65.8183
R4007 VGND.n2393 VGND.t86 65.8183
R4008 VGND.n2689 VGND.t80 65.8183
R4009 VGND.n2424 VGND.t86 65.8183
R4010 VGND.n2182 VGND.t86 65.8183
R4011 VGND.n2209 VGND.t86 65.8183
R4012 VGND.n2212 VGND.t86 65.8183
R4013 VGND.n2133 VGND.t80 65.8183
R4014 VGND.n2202 VGND.t80 65.8183
R4015 VGND.n2204 VGND.t80 65.8183
R4016 VGND.n2431 VGND.t80 65.8183
R4017 VGND.n1946 VGND.t81 65.8183
R4018 VGND.n1614 VGND.t81 65.8183
R4019 VGND.n1958 VGND.t81 65.8183
R4020 VGND.n1971 VGND.t81 65.8183
R4021 VGND.n1984 VGND.t81 65.8183
R4022 VGND.n1986 VGND.t81 65.8183
R4023 VGND.n2002 VGND.t81 65.8183
R4024 VGND.n2022 VGND.t81 65.8183
R4025 VGND.n2036 VGND.t81 65.8183
R4026 VGND.n2046 VGND.t81 65.8183
R4027 VGND.n2056 VGND.t81 65.8183
R4028 VGND.t83 VGND.n2327 65.8183
R4029 VGND.t83 VGND.n1053 65.8183
R4030 VGND.t83 VGND.n1052 65.8183
R4031 VGND.t83 VGND.n1051 65.8183
R4032 VGND.n2087 VGND.t77 65.8183
R4033 VGND.n2093 VGND.t77 65.8183
R4034 VGND.n2095 VGND.t77 65.8183
R4035 VGND.t83 VGND.n1042 65.8183
R4036 VGND.t83 VGND.n1049 65.8183
R4037 VGND.t83 VGND.n1040 65.8183
R4038 VGND.t83 VGND.n1050 65.8183
R4039 VGND.t83 VGND.n1048 65.8183
R4040 VGND.t83 VGND.n1047 65.8183
R4041 VGND.t83 VGND.n1046 65.8183
R4042 VGND.t83 VGND.n1045 65.8183
R4043 VGND.n2105 VGND.t77 65.8183
R4044 VGND.n2280 VGND.t77 65.8183
R4045 VGND.n2128 VGND.t77 65.8183
R4046 VGND.n2266 VGND.t77 65.8183
R4047 VGND.n2156 VGND.t77 65.8183
R4048 VGND.n2802 VGND.t77 65.8183
R4049 VGND.n518 VGND.t77 65.8183
R4050 VGND.n2843 VGND.t77 65.8183
R4051 VGND.n2838 VGND.t85 65.8183
R4052 VGND.n505 VGND.t85 65.8183
R4053 VGND.n2797 VGND.t85 65.8183
R4054 VGND.n523 VGND.t85 65.8183
R4055 VGND.n2452 VGND.t80 65.8183
R4056 VGND.n2467 VGND.t80 65.8183
R4057 VGND.n2764 VGND.t80 65.8183
R4058 VGND.t80 VGND.n575 65.8183
R4059 VGND.t79 VGND.n2774 65.8183
R4060 VGND.t79 VGND.n564 65.8183
R4061 VGND.t79 VGND.n563 65.8183
R4062 VGND.t79 VGND.n562 65.8183
R4063 VGND.n2229 VGND.t86 65.8183
R4064 VGND.n1037 VGND.t86 65.8183
R4065 VGND.n2338 VGND.t86 65.8183
R4066 VGND.n2335 VGND.t86 65.8183
R4067 VGND.n2734 VGND.t80 65.8183
R4068 VGND.n2173 VGND.t80 65.8183
R4069 VGND.n2171 VGND.t80 65.8183
R4070 VGND.n2259 VGND.t80 65.8183
R4071 VGND.t79 VGND.n554 65.8183
R4072 VGND.t79 VGND.n552 65.8183
R4073 VGND.t79 VGND.n550 65.8183
R4074 VGND.n2775 VGND.t79 65.8183
R4075 VGND.t83 VGND.n1043 65.8183
R4076 VGND.t83 VGND.n1041 65.8183
R4077 VGND.n2330 VGND.t83 65.8183
R4078 VGND.t83 VGND.n1029 65.8183
R4079 VGND.n2161 VGND.t77 65.8183
R4080 VGND.n2164 VGND.t77 65.8183
R4081 VGND.n2167 VGND.t77 65.8183
R4082 VGND.n2154 VGND.t77 65.8183
R4083 VGND.n651 VGND.t85 65.8183
R4084 VGND.n649 VGND.t85 65.8183
R4085 VGND.n627 VGND.t85 65.8183
R4086 VGND.n625 VGND.t85 65.8183
R4087 VGND.n2887 VGND.t81 65.8183
R4088 VGND.n464 VGND.t81 65.8183
R4089 VGND.n2904 VGND.t81 65.8183
R4090 VGND.t81 VGND.n441 65.8183
R4091 VGND.t84 VGND.n429 65.8183
R4092 VGND.t84 VGND.n428 65.8183
R4093 VGND.t84 VGND.n427 65.8183
R4094 VGND.t84 VGND.n426 65.8183
R4095 VGND.n90 VGND.n55 65.6721
R4096 VGND.n1463 VGND.n1462 65.4164
R4097 VGND.n2591 VGND.n951 65.3108
R4098 VGND.n3106 VGND.n194 65.0967
R4099 VGND.n114 VGND.n94 65.0005
R4100 VGND.n94 VGND.t42 65.0005
R4101 VGND.n101 VGND.n95 65.0005
R4102 VGND.n95 VGND.t42 65.0005
R4103 VGND.n98 VGND.n96 65.0005
R4104 VGND.n98 VGND.t118 65.0005
R4105 VGND.n107 VGND.n106 65.0005
R4106 VGND.n107 VGND.t118 65.0005
R4107 VGND.n946 VGND.n782 64.5959
R4108 VGND.t79 VGND.n557 64.1729
R4109 VGND.n2963 VGND.t85 64.1729
R4110 VGND.n1468 VGND.n1377 63.9439
R4111 VGND.n1565 VGND.n1564 61.901
R4112 VGND.n138 VGND.n123 61.6951
R4113 VGND.t78 VGND.n381 61.4728
R4114 VGND.t78 VGND.n2932 61.4728
R4115 VGND.n1255 VGND.n1254 61.1327
R4116 VGND.t14 VGND.t55 60.9543
R4117 VGND.n1206 VGND.n1178 60.4258
R4118 VGND.n115 VGND.n114 58.9497
R4119 VGND.n1193 VGND.n1179 58.6609
R4120 VGND.n2391 VGND.t86 57.8461
R4121 VGND.n2433 VGND.t80 57.8461
R4122 VGND.t79 VGND.n561 57.8461
R4123 VGND.t83 VGND.n1028 57.8461
R4124 VGND.n3283 VGND.n3282 56.6982
R4125 VGND.n2963 VGND.n2962 56.6572
R4126 VGND.n2964 VGND.n2963 56.6572
R4127 VGND.n2516 VGND.n557 56.6572
R4128 VGND.t95 VGND.n3106 56.5841
R4129 VGND.n1995 VGND.n1994 56.3995
R4130 VGND.n2714 VGND.n688 56.3995
R4131 VGND.n1994 VGND.n1066 56.3995
R4132 VGND.n1571 VGND.n1003 56.3995
R4133 VGND.n2554 VGND.n2553 56.3995
R4134 VGND.n2547 VGND.n2546 56.3995
R4135 VGND.n2936 VGND.n2935 56.3995
R4136 VGND.n2440 VGND.n2439 56.3995
R4137 VGND.n2700 VGND.n703 56.3995
R4138 VGND.n590 VGND.n589 56.3995
R4139 VGND.n591 VGND.n590 56.3995
R4140 VGND.n2721 VGND.n2720 56.3995
R4141 VGND.n541 VGND.n536 56.3995
R4142 VGND.n1572 VGND.n1571 56.3995
R4143 VGND.n1712 VGND.n1023 56.3995
R4144 VGND.n1185 VGND.n1184 56.2807
R4145 VGND.t114 VGND.n1436 56.1284
R4146 VGND.t123 VGND.n1436 56.1284
R4147 VGND.n1529 VGND.n1318 55.7181
R4148 VGND.n1529 VGND.n1528 55.7181
R4149 VGND.n1528 VGND.n1319 55.7181
R4150 VGND.n1323 VGND.n1319 55.7181
R4151 VGND.n1372 VGND.n1323 55.7181
R4152 VGND.n1372 VGND.n1344 55.7181
R4153 VGND.n1516 VGND.n1344 55.7181
R4154 VGND.n1516 VGND.n1515 55.7181
R4155 VGND.n1515 VGND.n1345 55.7181
R4156 VGND.n1349 VGND.n1345 55.7181
R4157 VGND.n1506 VGND.n1349 55.7181
R4158 VGND.n1506 VGND.n1505 55.7181
R4159 VGND.n1505 VGND.n1363 55.7181
R4160 VGND.n1364 VGND.n1363 55.7181
R4161 VGND.n1119 VGND.n1118 55.7181
R4162 VGND.n1132 VGND.n1118 55.7181
R4163 VGND.n1133 VGND.n1132 55.7181
R4164 VGND.n1134 VGND.n1133 55.7181
R4165 VGND.n1134 VGND.n1101 55.7181
R4166 VGND.n1142 VGND.n1101 55.7181
R4167 VGND.n1143 VGND.n1142 55.7181
R4168 VGND.n1144 VGND.n1143 55.7181
R4169 VGND.n1144 VGND.n258 55.7181
R4170 VGND.n3048 VGND.n258 55.7181
R4171 VGND.n3049 VGND.n3048 55.7181
R4172 VGND.n3050 VGND.n3049 55.7181
R4173 VGND.n3050 VGND.n240 55.7181
R4174 VGND.n3058 VGND.n240 55.7181
R4175 VGND.n3059 VGND.n3058 55.7181
R4176 VGND.n3060 VGND.n3059 55.7181
R4177 VGND.n3060 VGND.n225 55.7181
R4178 VGND.n3074 VGND.n225 55.7181
R4179 VGND.t84 VGND.n412 55.2026
R4180 VGND.t82 VGND.n287 55.2026
R4181 VGND.n2085 VGND.t77 55.2026
R4182 VGND.t83 VGND.n1044 55.2026
R4183 VGND.n2253 VGND.t86 55.2026
R4184 VGND.n599 VGND.t80 55.2026
R4185 VGND.n1624 VGND.t81 55.2026
R4186 VGND.n131 VGND.n129 54.9635
R4187 VGND.n143 VGND.n142 54.9635
R4188 VGND.n1895 VGND.t82 54.4705
R4189 VGND.n1082 VGND.t81 54.4705
R4190 VGND.n2102 VGND.t77 54.4705
R4191 VGND.n2835 VGND.t85 54.4705
R4192 VGND.t84 VGND.n2915 54.4705
R4193 VGND.n3261 VGND.n3260 54.1447
R4194 VGND.n65 VGND.n58 53.6894
R4195 VGND.n2313 VGND.n1050 53.3664
R4196 VGND.n2310 VGND.n1040 53.3664
R4197 VGND.n2306 VGND.n1049 53.3664
R4198 VGND.n2302 VGND.n1042 53.3664
R4199 VGND.n2286 VGND.n1045 53.3664
R4200 VGND.n2113 VGND.n1046 53.3664
R4201 VGND.n2271 VGND.n1047 53.3664
R4202 VGND.n2248 VGND.n1048 53.3664
R4203 VGND.n2347 VGND.n1029 53.3664
R4204 VGND.n2330 VGND.n2329 53.3664
R4205 VGND.n1041 VGND.n1039 53.3664
R4206 VGND.n2236 VGND.n1043 53.3664
R4207 VGND.n2327 VGND.n2326 53.3664
R4208 VGND.n1055 VGND.n1053 53.3664
R4209 VGND.n1732 VGND.n1052 53.3664
R4210 VGND.n1724 VGND.n1051 53.3664
R4211 VGND.n2335 VGND.n1015 53.3664
R4212 VGND.n2338 VGND.n2337 53.3664
R4213 VGND.n2334 VGND.n1037 53.3664
R4214 VGND.n2230 VGND.n2229 53.3664
R4215 VGND.n2212 VGND.n2211 53.3664
R4216 VGND.n2209 VGND.n2208 53.3664
R4217 VGND.n2182 VGND.n985 53.3664
R4218 VGND.n2424 VGND.n2423 53.3664
R4219 VGND.n2394 VGND.n2393 53.3664
R4220 VGND.n2406 VGND.n2405 53.3664
R4221 VGND.n2409 VGND.n2408 53.3664
R4222 VGND.n2421 VGND.n2420 53.3664
R4223 VGND.n2361 VGND.n2360 53.3664
R4224 VGND.n2363 VGND.n2362 53.3664
R4225 VGND.n2376 VGND.n2375 53.3664
R4226 VGND.n2379 VGND.n2378 53.3664
R4227 VGND.n2257 VGND.n2133 53.3664
R4228 VGND.n2202 VGND.n2201 53.3664
R4229 VGND.n2205 VGND.n2204 53.3664
R4230 VGND.n2431 VGND.n2430 53.3664
R4231 VGND.n2259 VGND.n2258 53.3664
R4232 VGND.n2171 VGND.n2132 53.3664
R4233 VGND.n2174 VGND.n2173 53.3664
R4234 VGND.n2734 VGND.n2733 53.3664
R4235 VGND.n2766 VGND.n575 53.3664
R4236 VGND.n2764 VGND.n2763 53.3664
R4237 VGND.n2474 VGND.n2467 53.3664
R4238 VGND.n2563 VGND.n2452 53.3664
R4239 VGND.n2690 VGND.n2689 53.3664
R4240 VGND.n2571 VGND.n713 53.3664
R4241 VGND.n2574 VGND.n2573 53.3664
R4242 VGND.n2561 VGND.n965 53.3664
R4243 VGND.n2776 VGND.n2775 53.3664
R4244 VGND.n635 VGND.n550 53.3664
R4245 VGND.n618 VGND.n552 53.3664
R4246 VGND.n656 VGND.n554 53.3664
R4247 VGND.n2774 VGND.n2773 53.3664
R4248 VGND.n573 VGND.n564 53.3664
R4249 VGND.n2760 VGND.n563 53.3664
R4250 VGND.n2468 VGND.n562 53.3664
R4251 VGND.n2538 VGND.n549 53.3664
R4252 VGND.n2533 VGND.n551 53.3664
R4253 VGND.n2497 VGND.n553 53.3664
R4254 VGND.n1886 VGND.n413 53.3664
R4255 VGND.n1772 VGND.n414 53.3664
R4256 VGND.n1872 VGND.n415 53.3664
R4257 VGND.n1789 VGND.n416 53.3664
R4258 VGND.n2918 VGND.n409 53.3664
R4259 VGND.n2916 VGND.n411 53.3664
R4260 VGND.n2861 VGND.n419 53.3664
R4261 VGND.n1788 VGND.n417 53.3664
R4262 VGND.n2860 VGND.n417 53.3664
R4263 VGND.n477 VGND.n419 53.3664
R4264 VGND.n2917 VGND.n2916 53.3664
R4265 VGND.n423 VGND.n409 53.3664
R4266 VGND.n431 VGND.n429 53.3664
R4267 VGND.n445 VGND.n428 53.3664
R4268 VGND.n2899 VGND.n427 53.3664
R4269 VGND.n462 VGND.n426 53.3664
R4270 VGND.n1921 VGND.n421 53.3664
R4271 VGND.n1646 VGND.n420 53.3664
R4272 VGND.n1910 VGND.n418 53.3664
R4273 VGND.n3022 VGND.n3021 53.3664
R4274 VGND.n827 VGND.n824 53.3664
R4275 VGND.n3013 VGND.n307 53.3664
R4276 VGND.n3011 VGND.n3010 53.3664
R4277 VGND.n1847 VGND.n1786 53.3664
R4278 VGND.n1837 VGND.n1805 53.3664
R4279 VGND.n1836 VGND.n1815 53.3664
R4280 VGND.n1828 VGND.n1827 53.3664
R4281 VGND.n1764 VGND.n1699 53.3664
R4282 VGND.n1882 VGND.n1881 53.3664
R4283 VGND.n1784 VGND.n1766 53.3664
R4284 VGND.n1868 VGND.n1867 53.3664
R4285 VGND.n1698 VGND.n1656 53.3664
R4286 VGND.n1687 VGND.n1686 53.3664
R4287 VGND.n1684 VGND.n1664 53.3664
R4288 VGND.n1672 VGND.n1664 53.3664
R4289 VGND.n1688 VGND.n1687 53.3664
R4290 VGND.n1685 VGND.n1656 53.3664
R4291 VGND.n1647 VGND.n418 53.3664
R4292 VGND.n1920 VGND.n420 53.3664
R4293 VGND.n1924 VGND.n421 53.3664
R4294 VGND.n1871 VGND.n416 53.3664
R4295 VGND.n1773 VGND.n415 53.3664
R4296 VGND.n1885 VGND.n414 53.3664
R4297 VGND.n1756 VGND.n413 53.3664
R4298 VGND.n1765 VGND.n1764 53.3664
R4299 VGND.n1881 VGND.n1880 53.3664
R4300 VGND.n1785 VGND.n1784 53.3664
R4301 VGND.n1867 VGND.n1866 53.3664
R4302 VGND.n1827 VGND.n309 53.3664
R4303 VGND.n1826 VGND.n1815 53.3664
R4304 VGND.n1838 VGND.n1837 53.3664
R4305 VGND.n1848 VGND.n1847 53.3664
R4306 VGND.n3012 VGND.n3011 53.3664
R4307 VGND.n826 VGND.n307 53.3664
R4308 VGND.n824 VGND.n289 53.3664
R4309 VGND.n3023 VGND.n3022 53.3664
R4310 VGND.n2508 VGND.n559 53.3664
R4311 VGND.n2986 VGND.n2985 53.3664
R4312 VGND.n337 VGND.n335 53.3664
R4313 VGND.n2974 VGND.n2973 53.3664
R4314 VGND.n347 VGND.n346 53.3664
R4315 VGND.n346 VGND.n338 53.3664
R4316 VGND.n2975 VGND.n2974 53.3664
R4317 VGND.n335 VGND.n326 53.3664
R4318 VGND.n2987 VGND.n2986 53.3664
R4319 VGND.n625 VGND.n624 53.3664
R4320 VGND.n628 VGND.n627 53.3664
R4321 VGND.n649 VGND.n648 53.3664
R4322 VGND.n652 VGND.n651 53.3664
R4323 VGND.n2838 VGND.n2837 53.3664
R4324 VGND.n2813 VGND.n505 53.3664
R4325 VGND.n2797 VGND.n2796 53.3664
R4326 VGND.n2794 VGND.n523 53.3664
R4327 VGND.n2828 VGND.n2814 53.3664
R4328 VGND.n2827 VGND.n2826 53.3664
R4329 VGND.n2820 VGND.n2816 53.3664
R4330 VGND.n2821 VGND.n2820 53.3664
R4331 VGND.n2826 VGND.n2825 53.3664
R4332 VGND.n2829 VGND.n2828 53.3664
R4333 VGND.n2562 VGND.n2561 53.3664
R4334 VGND.n2575 VGND.n2574 53.3664
R4335 VGND.n2572 VGND.n2571 53.3664
R4336 VGND.n2523 VGND.n553 53.3664
R4337 VGND.n2496 VGND.n551 53.3664
R4338 VGND.n2534 VGND.n549 53.3664
R4339 VGND.n2360 VGND.n2359 53.3664
R4340 VGND.n2362 VGND.n1008 53.3664
R4341 VGND.n2377 VGND.n2376 53.3664
R4342 VGND.n2378 VGND.n1000 53.3664
R4343 VGND.n2422 VGND.n2421 53.3664
R4344 VGND.n2408 VGND.n986 53.3664
R4345 VGND.n2407 VGND.n2406 53.3664
R4346 VGND.n2393 VGND.n993 53.3664
R4347 VGND.n2689 VGND.n2688 53.3664
R4348 VGND.n2425 VGND.n2424 53.3664
R4349 VGND.n2183 VGND.n2182 53.3664
R4350 VGND.n2210 VGND.n2209 53.3664
R4351 VGND.n2213 VGND.n2212 53.3664
R4352 VGND.n2198 VGND.n2133 53.3664
R4353 VGND.n2203 VGND.n2202 53.3664
R4354 VGND.n2204 VGND.n981 53.3664
R4355 VGND.n2432 VGND.n2431 53.3664
R4356 VGND.n2906 VGND.n441 53.3664
R4357 VGND.n2904 VGND.n2903 53.3664
R4358 VGND.n465 VGND.n464 53.3664
R4359 VGND.n2887 VGND.n2886 53.3664
R4360 VGND.n2057 VGND.n2056 53.3664
R4361 VGND.n2047 VGND.n2046 53.3664
R4362 VGND.n2036 VGND.n2013 53.3664
R4363 VGND.n2035 VGND.n2022 53.3664
R4364 VGND.n1972 VGND.n1971 53.3664
R4365 VGND.n1984 VGND.n1983 53.3664
R4366 VGND.n1987 VGND.n1986 53.3664
R4367 VGND.n2002 VGND.n2001 53.3664
R4368 VGND.n1959 VGND.n1958 53.3664
R4369 VGND.n1614 VGND.n1606 53.3664
R4370 VGND.n1947 VGND.n1946 53.3664
R4371 VGND.n1946 VGND.n1945 53.3664
R4372 VGND.n1615 VGND.n1614 53.3664
R4373 VGND.n1958 VGND.n1957 53.3664
R4374 VGND.n1971 VGND.n1076 53.3664
R4375 VGND.n1985 VGND.n1984 53.3664
R4376 VGND.n1986 VGND.n1071 53.3664
R4377 VGND.n2003 VGND.n2002 53.3664
R4378 VGND.n2022 VGND.n466 53.3664
R4379 VGND.n2037 VGND.n2036 53.3664
R4380 VGND.n2046 VGND.n2045 53.3664
R4381 VGND.n2056 VGND.n2055 53.3664
R4382 VGND.n2327 VGND.n1054 53.3664
R4383 VGND.n1733 VGND.n1053 53.3664
R4384 VGND.n1723 VGND.n1052 53.3664
R4385 VGND.n1720 VGND.n1051 53.3664
R4386 VGND.n2843 VGND.n2842 53.3664
R4387 VGND.n519 VGND.n518 53.3664
R4388 VGND.n2802 VGND.n2801 53.3664
R4389 VGND.n2157 VGND.n2156 53.3664
R4390 VGND.n2154 VGND.n2130 53.3664
R4391 VGND.n2168 VGND.n2167 53.3664
R4392 VGND.n2165 VGND.n2164 53.3664
R4393 VGND.n2162 VGND.n2161 53.3664
R4394 VGND.n2105 VGND.n2104 53.3664
R4395 VGND.n2281 VGND.n2280 53.3664
R4396 VGND.n2128 VGND.n2107 53.3664
R4397 VGND.n2267 VGND.n2266 53.3664
R4398 VGND.n2095 VGND.n2082 53.3664
R4399 VGND.n2094 VGND.n2093 53.3664
R4400 VGND.n2087 VGND.n2084 53.3664
R4401 VGND.n2088 VGND.n2087 53.3664
R4402 VGND.n2093 VGND.n2092 53.3664
R4403 VGND.n2096 VGND.n2095 53.3664
R4404 VGND.n2299 VGND.n1042 53.3664
R4405 VGND.n2303 VGND.n1049 53.3664
R4406 VGND.n2307 VGND.n1040 53.3664
R4407 VGND.n2311 VGND.n1050 53.3664
R4408 VGND.n2270 VGND.n1048 53.3664
R4409 VGND.n2114 VGND.n1047 53.3664
R4410 VGND.n2285 VGND.n1046 53.3664
R4411 VGND.n2074 VGND.n1045 53.3664
R4412 VGND.n2106 VGND.n2105 53.3664
R4413 VGND.n2280 VGND.n2279 53.3664
R4414 VGND.n2129 VGND.n2128 53.3664
R4415 VGND.n2266 VGND.n2265 53.3664
R4416 VGND.n2156 VGND.n520 53.3664
R4417 VGND.n2803 VGND.n2802 53.3664
R4418 VGND.n518 VGND.n502 53.3664
R4419 VGND.n2844 VGND.n2843 53.3664
R4420 VGND.n2839 VGND.n2838 53.3664
R4421 VGND.n2795 VGND.n505 53.3664
R4422 VGND.n2798 VGND.n2797 53.3664
R4423 VGND.n623 VGND.n523 53.3664
R4424 VGND.n2475 VGND.n2452 53.3664
R4425 VGND.n2467 VGND.n577 53.3664
R4426 VGND.n2765 VGND.n2764 53.3664
R4427 VGND.n597 VGND.n575 53.3664
R4428 VGND.n2774 VGND.n565 53.3664
R4429 VGND.n2759 VGND.n564 53.3664
R4430 VGND.n2469 VGND.n563 53.3664
R4431 VGND.n2465 VGND.n562 53.3664
R4432 VGND.n2229 VGND.n2214 53.3664
R4433 VGND.n2228 VGND.n1037 53.3664
R4434 VGND.n2339 VGND.n2338 53.3664
R4435 VGND.n2336 VGND.n2335 53.3664
R4436 VGND.n2735 VGND.n2734 53.3664
R4437 VGND.n2173 VGND.n601 53.3664
R4438 VGND.n2172 VGND.n2171 53.3664
R4439 VGND.n2260 VGND.n2259 53.3664
R4440 VGND.n2507 VGND.n554 53.3664
R4441 VGND.n655 VGND.n552 53.3664
R4442 VGND.n617 VGND.n550 53.3664
R4443 VGND.n2775 VGND.n548 53.3664
R4444 VGND.n2249 VGND.n1043 53.3664
R4445 VGND.n2235 VGND.n1041 53.3664
R4446 VGND.n2331 VGND.n2330 53.3664
R4447 VGND.n2328 VGND.n1029 53.3664
R4448 VGND.n2161 VGND.n2160 53.3664
R4449 VGND.n2164 VGND.n2163 53.3664
R4450 VGND.n2167 VGND.n2166 53.3664
R4451 VGND.n2155 VGND.n2154 53.3664
R4452 VGND.n651 VGND.n348 53.3664
R4453 VGND.n650 VGND.n649 53.3664
R4454 VGND.n627 VGND.n614 53.3664
R4455 VGND.n626 VGND.n625 53.3664
R4456 VGND.n2888 VGND.n2887 53.3664
R4457 VGND.n464 VGND.n443 53.3664
R4458 VGND.n2905 VGND.n2904 53.3664
R4459 VGND.n1622 VGND.n441 53.3664
R4460 VGND.n444 VGND.n429 53.3664
R4461 VGND.n2900 VGND.n428 53.3664
R4462 VGND.n461 VGND.n427 53.3664
R4463 VGND.n2883 VGND.n426 53.3664
R4464 VGND.n1389 VGND.n1377 51.2005
R4465 VGND.n2668 VGND.n728 50.7155
R4466 VGND.n1212 VGND.n1211 50.3571
R4467 VGND.n148 VGND.n147 50.3569
R4468 VGND.n1159 VGND.t10 50.3367
R4469 VGND.t21 VGND.n229 50.3367
R4470 VGND.n3189 VGND.n3154 49.9965
R4471 VGND.n2622 VGND.n2619 49.073
R4472 VGND.n3170 VGND.n3169 48.7507
R4473 VGND.n3186 VGND.n3185 48.7507
R4474 VGND.n2581 VGND.n956 48.7505
R4475 VGND.n2581 VGND.n2580 48.7505
R4476 VGND.n2586 VGND.n2585 48.7505
R4477 VGND.n2585 VGND.n947 48.7505
R4478 VGND.n2681 VGND.n2680 48.7505
R4479 VGND.n2682 VGND.n2681 48.7505
R4480 VGND.n1590 VGND.n1569 48.7505
R4481 VGND.n1598 VGND.n1569 48.7505
R4482 VGND.t50 VGND.t91 48.4465
R4483 VGND.t114 VGND.t69 48.4465
R4484 VGND.t34 VGND.t2 48.4465
R4485 VGND.t37 VGND.t103 48.4465
R4486 VGND.t59 VGND.t112 48.4465
R4487 VGND.t74 VGND.t105 48.4465
R4488 VGND.n101 VGND.n34 47.7763
R4489 VGND.n3210 VGND.n3209 47.4646
R4490 VGND.n3224 VGND.n3223 47.4646
R4491 VGND.n3215 VGND.n3214 47.4646
R4492 VGND.t9 VGND.n234 47.4265
R4493 VGND.t72 VGND.n1122 47.4265
R4494 VGND.t31 VGND.n1112 47.4265
R4495 VGND.t17 VGND.n1103 47.4265
R4496 VGND.t8 VGND.n1095 47.4265
R4497 VGND.t16 VGND.n260 47.4265
R4498 VGND.t12 VGND.n250 47.4265
R4499 VGND.t7 VGND.n242 47.4265
R4500 VGND.t21 VGND.n228 47.4265
R4501 VGND.n1122 VGND.t10 47.4265
R4502 VGND.t72 VGND.n1112 47.4265
R4503 VGND.t31 VGND.n1103 47.4265
R4504 VGND.t17 VGND.n1095 47.4265
R4505 VGND.t8 VGND.n260 47.4265
R4506 VGND.t16 VGND.n250 47.4265
R4507 VGND.t12 VGND.n242 47.4265
R4508 VGND.t9 VGND.n228 47.4265
R4509 VGND.n234 VGND.n221 46.4652
R4510 VGND.n1364 VGND.n12 46.3064
R4511 VGND.n1420 VGND.t57 46.3007
R4512 VGND.n3201 VGND.n3200 45.4342
R4513 VGND.t69 VGND.n1301 45.3808
R4514 VGND.n3200 VGND.n3154 44.8005
R4515 VGND.n829 VGND.t70 44.0166
R4516 VGND.n3210 VGND.n3147 43.9125
R4517 VGND.n3223 VGND.n83 43.9125
R4518 VGND.n3214 VGND.n48 43.9125
R4519 VGND.t57 VGND.n1404 43.5411
R4520 VGND.n3037 VGND.t71 43.3166
R4521 VGND.n3240 VGND.n48 43.3
R4522 VGND.n3169 VGND.n83 43.3
R4523 VGND.n3185 VGND.n3147 43.3
R4524 VGND.n152 VGND.n16 43.1245
R4525 VGND.n1458 VGND.n1318 42.9181
R4526 VGND.n1437 VGND.t114 42.6142
R4527 VGND.t123 VGND.n1437 42.6142
R4528 VGND.n829 VGND.t19 42.5516
R4529 VGND.n742 VGND.t101 42.5516
R4530 VGND.n740 VGND.t122 42.5516
R4531 VGND.n1595 VGND.n1580 42.51
R4532 VGND.n830 VGND.t18 42.3691
R4533 VGND.n739 VGND.t121 42.3691
R4534 VGND.n741 VGND.t100 42.3691
R4535 VGND.t58 VGND.n1300 42.3146
R4536 VGND.n1441 VGND.n1297 42.2536
R4537 VGND.n3035 VGND.n3034 41.9315
R4538 VGND.n2580 VGND.n2579 41.6984
R4539 VGND.n3284 VGND.n3283 41.3519
R4540 VGND.n1183 VGND.n1172 41.2394
R4541 VGND.n2515 VGND.n2514 41.2097
R4542 VGND.n1413 VGND.n1412 39.638
R4543 VGND.n1119 VGND.n1092 39.5299
R4544 VGND.n3075 VGND.n3074 39.5299
R4545 VGND.t104 VGND.n1294 39.2484
R4546 VGND.t103 VGND.n1397 39.2484
R4547 VGND.n2682 VGND.t78 39.0923
R4548 VGND.n1281 VGND.n1280 38.7219
R4549 VGND.t6 VGND.n759 38.5575
R4550 VGND.t78 VGND.n384 38.0567
R4551 VGND.n1444 VGND.n1405 37.976
R4552 VGND.n3264 VGND.n16 37.6559
R4553 VGND.n2669 VGND.n2668 37.3818
R4554 VGND.n960 VGND.t78 37.3549
R4555 VGND.n113 VGND.n96 37.1867
R4556 VGND.n114 VGND.n113 36.8557
R4557 VGND.n1438 VGND.t34 36.4888
R4558 VGND.n1255 VGND.n4 36.2511
R4559 VGND.t97 VGND.n1293 36.1822
R4560 VGND.n1256 VGND.n1255 35.8662
R4561 VGND.n1463 VGND.n1458 34.6624
R4562 VGND.n3168 VGND.n46 33.3552
R4563 VGND.t54 VGND.n1287 33.116
R4564 VGND.n3237 VGND.n58 32.5931
R4565 VGND.n966 VGND.n716 32.5005
R4566 VGND.n2682 VGND.n716 32.5005
R4567 VGND.n2598 VGND.n2597 32.5005
R4568 VGND.n2599 VGND.n2598 32.5005
R4569 VGND.n957 VGND.n720 32.5005
R4570 VGND.n958 VGND.n957 32.5005
R4571 VGND.n1597 VGND.n1596 32.5005
R4572 VGND.n1598 VGND.n1597 32.5005
R4573 VGND.n1213 VGND.n1163 32.5005
R4574 VGND.n1199 VGND.n1163 32.5005
R4575 VGND.n1268 VGND.n6 32.5005
R4576 VGND.n1269 VGND.n1268 32.5005
R4577 VGND.n1426 VGND.t59 32.1961
R4578 VGND.n2674 VGND.n2673 31.5562
R4579 VGND.n1078 VGND.n1062 31.4187
R4580 VGND.n1586 VGND.n956 31.1247
R4581 VGND.n67 VGND.n46 30.926
R4582 VGND.n3224 VGND.n82 30.5783
R4583 VGND.n2670 VGND.n725 30.4557
R4584 VGND.n960 VGND.n958 30.4052
R4585 VGND.n1192 VGND.n1191 30.188
R4586 VGND.t48 VGND.n1286 30.0498
R4587 VGND.n3215 VGND.n81 29.9857
R4588 VGND.n3209 VGND.n3149 29.6301
R4589 VGND.n3209 VGND.n3208 29.5116
R4590 VGND.n1458 VGND.n1457 29.5085
R4591 VGND.n3225 VGND.n3224 29.3931
R4592 VGND.n3185 VGND.n53 29.2505
R4593 VGND.t46 VGND.n53 29.2505
R4594 VGND.n3154 VGND.n54 29.2505
R4595 VGND.t46 VGND.n54 29.2505
R4596 VGND.n3210 VGND.n92 29.2505
R4597 VGND.t35 VGND.n92 29.2505
R4598 VGND.n3201 VGND.n93 29.2505
R4599 VGND.t35 VGND.n93 29.2505
R4600 VGND.n3169 VGND.n57 29.2505
R4601 VGND.t46 VGND.n57 29.2505
R4602 VGND.n3185 VGND.n56 29.2505
R4603 VGND.t46 VGND.n56 29.2505
R4604 VGND.n3223 VGND.n84 29.2505
R4605 VGND.t35 VGND.n84 29.2505
R4606 VGND.n3211 VGND.n3210 29.2505
R4607 VGND.t35 VGND.n3211 29.2505
R4608 VGND.n3240 VGND.n47 29.2505
R4609 VGND.t46 VGND.n47 29.2505
R4610 VGND.n3169 VGND.n52 29.2505
R4611 VGND.t46 VGND.n52 29.2505
R4612 VGND.n3214 VGND.n91 29.2505
R4613 VGND.t35 VGND.n91 29.2505
R4614 VGND.n3223 VGND.n3222 29.2505
R4615 VGND.n3222 VGND.t35 29.2505
R4616 VGND.n3238 VGND.n3237 29.2505
R4617 VGND.t46 VGND.n3238 29.2505
R4618 VGND.n3240 VGND.n3239 29.2505
R4619 VGND.n3239 VGND.t46 29.2505
R4620 VGND.n3221 VGND.n59 29.2505
R4621 VGND.t35 VGND.n3221 29.2505
R4622 VGND.n3214 VGND.n3212 29.2505
R4623 VGND.t35 VGND.n3212 29.2505
R4624 VGND.n2680 VGND.n719 29.1741
R4625 VGND.n1591 VGND.n1580 28.9016
R4626 VGND.n3218 VGND.n3215 28.3264
R4627 VGND.n137 VGND.n136 28.1893
R4628 VGND.n135 VGND.n24 28.1893
R4629 VGND.n139 VGND.n138 28.1893
R4630 VGND.n140 VGND.n137 28.1893
R4631 VGND.n140 VGND.n139 28.1893
R4632 VGND.n1564 VGND.n1273 28.1718
R4633 VGND.n136 VGND.n135 28.0454
R4634 VGND.n194 VGND.n188 28.0419
R4635 VGND.n66 VGND.n65 27.8428
R4636 VGND.n3241 VGND.n46 27.3766
R4637 VGND.n381 VGND.n353 27.1902
R4638 VGND.n2932 VGND.n316 27.1902
R4639 VGND.t62 VGND.n1278 26.9836
R4640 VGND.n1248 VGND.n1247 26.504
R4641 VGND.t126 VGND.n1161 25.8924
R4642 VGND.n106 VGND.n103 25.8304
R4643 VGND.n146 VGND.n145 25.6785
R4644 VGND.n103 VGND.n101 25.6005
R4645 VGND.n3266 VGND.n20 25.5229
R4646 VGND.t105 VGND.n1381 25.1439
R4647 VGND.n133 VGND.n29 24.9761
R4648 VGND.n1442 VGND.n1441 24.6209
R4649 VGND.n1277 VGND.t50 24.5306
R4650 VGND.t78 VGND.n380 24.4596
R4651 VGND.n3170 VGND.n3166 24.1056
R4652 VGND.t53 VGND.n1277 23.9174
R4653 VGND.n1247 VGND.n1185 23.5153
R4654 VGND.n3188 VGND.n3186 23.3582
R4655 VGND.t125 VGND.n1381 23.3041
R4656 VGND.n3186 VGND.n3184 23.2647
R4657 VGND.n3171 VGND.n3170 23.1713
R4658 VGND.n3283 VGND.n5 22.9687
R4659 VGND.n1213 VGND.n1212 22.6545
R4660 VGND.n1217 VGND.n1186 22.57
R4661 VGND.n3190 VGND.n3189 22.3068
R4662 VGND.n135 VGND.n19 21.7217
R4663 VGND.n139 VGND.n127 21.6981
R4664 VGND.n137 VGND.n28 21.542
R4665 VGND.n1278 VGND.t53 21.4644
R4666 VGND.n2933 VGND.t78 20.8495
R4667 VGND.n2674 VGND.n720 20.2726
R4668 VGND.n1203 VGND.n1202 20.1729
R4669 VGND.n1202 VGND.n1160 20.1729
R4670 VGND.n1196 VGND.n1188 20.1729
R4671 VGND.n1200 VGND.n1196 20.1729
R4672 VGND.n1197 VGND.n1185 20.1729
R4673 VGND.n1198 VGND.n1197 20.1729
R4674 VGND.n1167 VGND.n4 20.1729
R4675 VGND.n1167 VGND.n1161 20.1729
R4676 VGND.n1172 VGND.n1170 20.1729
R4677 VGND.n1198 VGND.n1170 20.1729
R4678 VGND.n1257 VGND.n1171 20.1729
R4679 VGND.n1171 VGND.n1161 20.1729
R4680 VGND.n1277 VGND.n1275 20.0282
R4681 VGND.n3176 VGND.n3147 19.9729
R4682 VGND.n1226 VGND.t39 19.8367
R4683 VGND.n1231 VGND.t127 19.8235
R4684 VGND.n3177 VGND.n3176 19.7522
R4685 VGND.n87 VGND.n83 19.5315
R4686 VGND.n1286 VGND.n1285 19.4978
R4687 VGND.n1254 VGND.n1176 19.4453
R4688 VGND.n3269 VGND.n3268 19.0262
R4689 VGND.n3162 VGND.n3157 18.9246
R4690 VGND.n3200 VGND.n3157 18.8143
R4691 VGND.n1286 VGND.t62 18.3982
R4692 VGND.n1441 VGND.n1440 18.2817
R4693 VGND.n1440 VGND.n1439 18.2817
R4694 VGND.n1424 VGND.n1423 18.2817
R4695 VGND.n1423 VGND.n1422 18.2817
R4696 VGND.n1430 VGND.n1429 18.2817
R4697 VGND.n1429 VGND.n1428 18.2817
R4698 VGND.n1380 VGND.n1377 18.2817
R4699 VGND.n1459 VGND.n1380 18.2817
R4700 VGND.n1405 VGND.n1401 18.2817
R4701 VGND.n1439 VGND.n1401 18.2817
R4702 VGND.n1421 VGND.n1399 18.2817
R4703 VGND.n1422 VGND.n1421 18.2817
R4704 VGND.n1427 VGND.n1391 18.2817
R4705 VGND.n1428 VGND.n1427 18.2817
R4706 VGND.n1457 VGND.n1385 18.2817
R4707 VGND.n1459 VGND.n1385 18.2817
R4708 VGND.n1293 VGND.n1292 17.7887
R4709 VGND.n1195 VGND.n1194 17.7278
R4710 VGND.t124 VGND.n1195 17.7278
R4711 VGND.n1201 VGND.n1190 17.7278
R4712 VGND.n1201 VGND.t124 17.7278
R4713 VGND.n1566 VGND.n1565 17.7278
R4714 VGND.n1567 VGND.n1566 17.7278
R4715 VGND.n1462 VGND.n1461 17.7278
R4716 VGND.n1461 VGND.n1460 17.7278
R4717 VGND.n1176 VGND.n1166 17.7278
R4718 VGND.t14 VGND.n1166 17.7278
R4719 VGND.n1168 VGND.n5 17.7278
R4720 VGND.t14 VGND.n1168 17.7278
R4721 VGND.n1265 VGND.n1264 17.7278
R4722 VGND.t14 VGND.n1265 17.7278
R4723 VGND.n1176 VGND.n1169 17.7278
R4724 VGND.t14 VGND.n1169 17.7278
R4725 VGND.n87 VGND.n85 17.5453
R4726 VGND.n3241 VGND.n3240 17.2101
R4727 VGND.n2504 VGND.n364 17.1825
R4728 VGND.n2509 VGND.n365 17.1825
R4729 VGND.n2597 VGND.n727 17.0672
R4730 VGND.n1464 VGND.n1463 16.6548
R4731 VGND.n1228 VGND.n1222 16.5104
R4732 VGND.n1227 VGND.n1224 16.5104
R4733 VGND.n1229 VGND.n1221 16.51
R4734 VGND.n968 VGND.n966 16.5058
R4735 VGND.n1232 VGND.n1230 16.4747
R4736 VGND.n62 VGND.n61 16.3867
R4737 VGND.n1426 VGND.t74 16.2519
R4738 VGND.n2832 VGND.n492 16.0005
R4739 VGND.n2832 VGND.n2831 16.0005
R4740 VGND.n2831 VGND.n2830 16.0005
R4741 VGND.n2830 VGND.n2815 16.0005
R4742 VGND.n2824 VGND.n2815 16.0005
R4743 VGND.n2824 VGND.n2823 16.0005
R4744 VGND.n2823 VGND.n2822 16.0005
R4745 VGND.n2822 VGND.n2819 16.0005
R4746 VGND.n2099 VGND.n2065 16.0005
R4747 VGND.n2099 VGND.n2098 16.0005
R4748 VGND.n2098 VGND.n2097 16.0005
R4749 VGND.n2097 VGND.n2083 16.0005
R4750 VGND.n2091 VGND.n2083 16.0005
R4751 VGND.n2091 VGND.n2090 16.0005
R4752 VGND.n2090 VGND.n2089 16.0005
R4753 VGND.n2089 VGND.n493 16.0005
R4754 VGND.n2314 VGND.n2312 16.0005
R4755 VGND.n2312 VGND.n2309 16.0005
R4756 VGND.n2309 VGND.n2308 16.0005
R4757 VGND.n2308 VGND.n2305 16.0005
R4758 VGND.n2305 VGND.n2304 16.0005
R4759 VGND.n2304 VGND.n2301 16.0005
R4760 VGND.n2301 VGND.n2300 16.0005
R4761 VGND.n2300 VGND.n2297 16.0005
R4762 VGND.n858 VGND.n779 15.8046
R4763 VGND.n3260 VGND.n20 15.6805
R4764 VGND.n126 VGND.n125 15.6805
R4765 VGND.n146 VGND.n126 15.6805
R4766 VGND.n125 VGND.n124 15.6805
R4767 VGND.n147 VGND.n146 15.6805
R4768 VGND.n124 VGND.n20 15.6005
R4769 VGND.n1287 VGND.t48 15.332
R4770 VGND.n2592 VGND.n2591 15.2016
R4771 VGND.n1300 VGND.n1299 14.9009
R4772 VGND.n2596 VGND.n950 14.8567
R4773 VGND.n1390 VGND.n1389 14.6695
R4774 VGND.n1217 VGND.n1162 14.6255
R4775 VGND.n1266 VGND.n1162 14.6255
R4776 VGND.n1267 VGND.n1165 14.6255
R4777 VGND.n1267 VGND.n1266 14.6255
R4778 VGND.n1448 VGND.n1400 14.57
R4779 VGND.n1184 VGND.n1183 14.5437
R4780 VGND.n3235 VGND.n62 14.5108
R4781 VGND.n838 VGND.n797 14.2688
R4782 VGND.t1 VGND.n838 14.2688
R4783 VGND.n2601 VGND.n2600 14.2688
R4784 VGND.n2600 VGND.t1 14.2688
R4785 VGND.n839 VGND.n810 14.2688
R4786 VGND.t1 VGND.n839 14.2688
R4787 VGND.n841 VGND.n314 14.2688
R4788 VGND.t1 VGND.n841 14.2688
R4789 VGND.n885 VGND.n843 14.2688
R4790 VGND.t1 VGND.n843 14.2688
R4791 VGND.n883 VGND.n845 14.2688
R4792 VGND.t1 VGND.n845 14.2688
R4793 VGND.n882 VGND.n847 14.2688
R4794 VGND.t1 VGND.n847 14.2688
R4795 VGND.n879 VGND.n849 14.2688
R4796 VGND.t1 VGND.n849 14.2688
R4797 VGND.n866 VGND.n851 14.2688
R4798 VGND.t1 VGND.n851 14.2688
R4799 VGND.n853 VGND.n366 14.2688
R4800 VGND.t1 VGND.n853 14.2688
R4801 VGND.n855 VGND.n363 14.2688
R4802 VGND.t1 VGND.n855 14.2688
R4803 VGND.n2615 VGND.n2614 14.2688
R4804 VGND.n2614 VGND.t6 14.2688
R4805 VGND.n836 VGND.n804 14.2688
R4806 VGND.n836 VGND.t6 14.2688
R4807 VGND.n2606 VGND.n2605 14.2688
R4808 VGND.n2606 VGND.t6 14.2688
R4809 VGND.n906 VGND.n905 14.2688
R4810 VGND.n905 VGND.t6 14.2688
R4811 VGND.n891 VGND.n886 14.2688
R4812 VGND.n891 VGND.t6 14.2688
R4813 VGND.n897 VGND.n884 14.2688
R4814 VGND.n897 VGND.t6 14.2688
R4815 VGND.n915 VGND.n914 14.2688
R4816 VGND.n915 VGND.t6 14.2688
R4817 VGND.n918 VGND.n869 14.2688
R4818 VGND.n918 VGND.t6 14.2688
R4819 VGND.n926 VGND.n925 14.2688
R4820 VGND.n926 VGND.t6 14.2688
R4821 VGND.n931 VGND.n930 14.2688
R4822 VGND.n930 VGND.t6 14.2688
R4823 VGND.n936 VGND.n935 14.2688
R4824 VGND.n936 VGND.t6 14.2688
R4825 VGND.n952 VGND.n945 14.2688
R4826 VGND.t1 VGND.n945 14.2688
R4827 VGND.n943 VGND.n942 14.2688
R4828 VGND.n943 VGND.t6 14.2688
R4829 VGND.n3034 VGND.n3033 14.2688
R4830 VGND.n3033 VGND.n3032 14.2688
R4831 VGND.n800 VGND.n799 14.2688
R4832 VGND.n799 VGND.n195 14.2688
R4833 VGND.n2623 VGND.n728 13.9485
R4834 VGND.n2623 VGND.n2621 13.9485
R4835 VGND.n2621 VGND.n767 13.9485
R4836 VGND.n2650 VGND.n767 13.9485
R4837 VGND.n2651 VGND.n2650 13.9485
R4838 VGND.n2652 VGND.n2651 13.9485
R4839 VGND.n2652 VGND.n757 13.9485
R4840 VGND.n2658 VGND.n757 13.9485
R4841 VGND.n2659 VGND.n2658 13.9485
R4842 VGND.n3118 VGND.n3117 13.9485
R4843 VGND.n3117 VGND.n3116 13.9485
R4844 VGND.n3116 VGND.n186 13.9485
R4845 VGND.n3107 VGND.n186 13.9485
R4846 VGND.n3107 VGND.n158 13.9485
R4847 VGND.n3137 VGND.n158 13.9485
R4848 VGND.n3138 VGND.n3137 13.9485
R4849 VGND.n3139 VGND.n3138 13.9485
R4850 VGND.n1449 VGND.n1448 13.9425
R4851 VGND.n1450 VGND.n1449 13.9425
R4852 VGND.n1450 VGND.n1386 13.9425
R4853 VGND.n1464 VGND.n1386 13.9425
R4854 VGND.n1214 VGND.n1188 13.918
R4855 VGND.n2317 VGND.n2316 13.8005
R4856 VGND.n70 VGND.n65 13.7852
R4857 VGND.n881 VGND.n880 13.7148
R4858 VGND.n2617 VGND.n277 13.7148
R4859 VGND.n1535 VGND.n1534 13.6533
R4860 VGND.n1468 VGND.n1467 13.6175
R4861 VGND.n1536 VGND.n1535 13.6091
R4862 VGND.n2617 VGND.n2616 13.5842
R4863 VGND.n966 VGND.n956 13.4742
R4864 VGND.n861 VGND.n859 13.4536
R4865 VGND.n1443 VGND.n1442 13.3556
R4866 VGND.n2602 VGND.n795 13.1923
R4867 VGND.n103 VGND.n102 12.9706
R4868 VGND.n2604 VGND.n2603 12.9311
R4869 VGND.n1188 VGND.n1186 12.8921
R4870 VGND.n922 VGND.n921 12.8805
R4871 VGND.n801 VGND.n798 12.8005
R4872 VGND.n934 VGND.n933 12.7205
R4873 VGND.n113 VGND.n112 12.6304
R4874 VGND.n2611 VGND.n2610 12.5605
R4875 VGND.n907 VGND.n808 12.5393
R4876 VGND.n873 VGND.n868 12.4087
R4877 VGND.n912 VGND.n911 12.4087
R4878 VGND.n2609 VGND.n805 12.4005
R4879 VGND.n913 VGND.n912 12.2781
R4880 VGND.n1293 VGND.t54 12.2658
R4881 VGND.n953 VGND.n952 12.1878
R4882 VGND.n888 VGND.n887 12.1605
R4883 VGND.n909 VGND.n908 12.1474
R4884 VGND.n862 VGND.n861 12.1474
R4885 VGND.n924 VGND.n923 12.0805
R4886 VGND.n910 VGND.n909 12.0168
R4887 VGND.n867 VGND.n862 12.0168
R4888 VGND.n893 VGND.n870 12.0005
R4889 VGND.n1438 VGND.t123 11.9592
R4890 VGND.n902 VGND.n901 11.9205
R4891 VGND.n913 VGND.n881 11.8862
R4892 VGND.n932 VGND.n860 11.8405
R4893 VGND.n933 VGND.n932 11.8405
R4894 VGND.n901 VGND.n900 11.7605
R4895 VGND.n911 VGND.n910 11.7556
R4896 VGND.n868 VGND.n867 11.7556
R4897 VGND.n900 VGND.n895 11.6805
R4898 VGND.n921 VGND.n870 11.6805
R4899 VGND.n908 VGND.n907 11.625
R4900 VGND.n2586 VGND.n778 11.6226
R4901 VGND.n924 VGND.n860 11.6005
R4902 VGND.n1412 VGND.n1281 11.5512
R4903 VGND.n902 VGND.n888 11.5205
R4904 VGND.n1417 VGND.n1406 11.3999
R4905 VGND.n1417 VGND.n1416 11.3999
R4906 VGND.n1467 VGND.n1378 11.3999
R4907 VGND.n1416 VGND.n1415 11.3221
R4908 VGND.n887 VGND.n805 11.2805
R4909 VGND.n380 VGND.n283 11.2426
R4910 VGND.n2604 VGND.n808 11.2332
R4911 VGND.n2610 VGND.n2609 11.1205
R4912 VGND.n1536 VGND.n1270 11.0382
R4913 VGND.n1436 VGND.n1270 11.0382
R4914 VGND.n1400 VGND.n1271 11.0382
R4915 VGND.n1437 VGND.n1271 11.0382
R4916 VGND.n2680 VGND.n2679 10.9812
R4917 VGND.n2603 VGND.n2602 10.9719
R4918 VGND.n934 VGND.n190 10.9605
R4919 VGND.n2611 VGND.n798 10.8805
R4920 VGND.n1292 VGND.n1289 10.8338
R4921 VGND.n1285 VGND.n1282 10.8338
R4922 VGND.n1442 VGND.n1298 10.8338
R4923 VGND.t69 VGND.n1298 10.8338
R4924 VGND.n1299 VGND.n1296 10.8338
R4925 VGND.n1280 VGND.n1275 10.8338
R4926 VGND.n1588 VGND.n1587 10.8149
R4927 VGND.n923 VGND.n922 10.8005
R4928 VGND.n1406 VGND.n1297 10.7385
R4929 VGND.n859 VGND.n858 10.7107
R4930 VGND.n2616 VGND.n795 10.5801
R4931 VGND.n880 VGND.n873 10.4495
R4932 VGND.n3112 VGND.n190 10.1605
R4933 VGND.n2583 VGND.n951 10.0718
R4934 VGND.n2851 VGND.n493 9.95606
R4935 VGND.n2297 VGND.n2296 9.95606
R4936 VGND.n1497 VGND.n1496 9.91575
R4937 VGND.n1496 VGND.n23 9.91575
R4938 VGND.n1501 VGND.n1500 9.91575
R4939 VGND.n1501 VGND.n1494 9.91575
R4940 VGND.n1508 VGND.n1507 9.91575
R4941 VGND.n1507 VGND.n1354 9.91575
R4942 VGND.n1357 VGND.n1347 9.91575
R4943 VGND.n1350 VGND.n1347 9.91575
R4944 VGND.n1518 VGND.n1517 9.91575
R4945 VGND.n1519 VGND.n1518 9.91575
R4946 VGND.n1336 VGND.n1335 9.91575
R4947 VGND.n1335 VGND.n1328 9.91575
R4948 VGND.n1331 VGND.n1321 9.91575
R4949 VGND.n1324 VGND.n1321 9.91575
R4950 VGND.n1531 VGND.n1530 9.91575
R4951 VGND.n1532 VGND.n1531 9.91575
R4952 VGND.n1309 VGND.n1307 9.91575
R4953 VGND.n1311 VGND.n1309 9.91575
R4954 VGND.n1490 VGND.n1489 9.91575
R4955 VGND.n1489 VGND.n1367 9.91575
R4956 VGND.n1368 VGND.n1362 9.91575
R4957 VGND.n1368 VGND.n1351 9.91575
R4958 VGND.n1371 VGND.n1346 9.91575
R4959 VGND.n1353 VGND.n1346 9.91575
R4960 VGND.n1481 VGND.n1343 9.91575
R4961 VGND.n1481 VGND.n1339 9.91575
R4962 VGND.n1375 VGND.n1374 9.91575
R4963 VGND.n1374 VGND.n1325 9.91575
R4964 VGND.n1376 VGND.n1320 9.91575
R4965 VGND.n1327 VGND.n1320 9.91575
R4966 VGND.n1471 VGND.n1317 9.91575
R4967 VGND.n1471 VGND.n1312 9.91575
R4968 VGND.n3272 VGND.n3271 9.91575
R4969 VGND.n3271 VGND.n3270 9.91575
R4970 VGND.n1389 VGND.n1388 9.91575
R4971 VGND.n1388 VGND.n1315 9.91575
R4972 VGND.n2951 VGND.n364 9.8023
R4973 VGND.n2951 VGND.n365 9.8023
R4974 VGND.n2506 VGND.n359 9.73111
R4975 VGND.n1247 VGND.n1246 9.59552
R4976 VGND.n955 VGND.n360 9.59066
R4977 VGND.n955 VGND.t107 9.59066
R4978 VGND.n766 VGND.n765 9.59066
R4979 VGND.n765 VGND.n763 9.59066
R4980 VGND.n939 VGND.n760 9.59066
R4981 VGND.n760 VGND.n759 9.59066
R4982 VGND.n756 VGND.n755 9.59066
R4983 VGND.n755 VGND.n179 9.59066
R4984 VGND.n185 VGND.n184 9.59066
R4985 VGND.n184 VGND.n180 9.59066
R4986 VGND.n746 VGND.n745 9.59066
R4987 VGND.n745 VGND.n161 9.59066
R4988 VGND.n772 VGND.n771 9.59066
R4989 VGND.n771 VGND.n769 9.59066
R4990 VGND.n2624 VGND.n2620 9.59066
R4991 VGND.n2622 VGND.n2620 9.59066
R4992 VGND.n3141 VGND.n3140 9.59066
R4993 VGND.n3142 VGND.n3141 9.59066
R4994 VGND.n193 VGND.n192 9.59066
R4995 VGND.n194 VGND.n193 9.59066
R4996 VGND.n164 VGND.n157 9.59066
R4997 VGND.n164 VGND.n162 9.59066
R4998 VGND.n950 VGND.n780 9.59066
R4999 VGND.n782 VGND.n780 9.59066
R5000 VGND.n949 VGND.n725 9.59066
R5001 VGND.n949 VGND.t52 9.59066
R5002 VGND.n2582 VGND.n948 9.59066
R5003 VGND.t52 VGND.n948 9.59066
R5004 VGND.n2584 VGND.n2583 9.59066
R5005 VGND.n2584 VGND.t107 9.59066
R5006 VGND.n1587 VGND.n717 9.59066
R5007 VGND.t22 VGND.n717 9.59066
R5008 VGND.n1589 VGND.n718 9.59066
R5009 VGND.t22 VGND.n718 9.59066
R5010 VGND.n1582 VGND.n1577 9.59066
R5011 VGND.n1577 VGND.t22 9.59066
R5012 VGND.n1587 VGND.n1578 9.59066
R5013 VGND.n1578 VGND.t22 9.59066
R5014 VGND.n273 VGND.n272 9.54799
R5015 VGND.n272 VGND.t133 9.53872
R5016 VGND.n271 VGND.t131 9.53872
R5017 VGND.n2502 VGND.n362 9.39557
R5018 VGND.n2588 VGND.n778 9.37714
R5019 VGND.n30 VGND 9.35119
R5020 VGND.n1154 VGND.n209 9.3005
R5021 VGND.n1149 VGND.n1148 9.3005
R5022 VGND.n2676 VGND.n2675 9.3005
R5023 VGND.n3189 VGND.n3158 9.3005
R5024 VGND.n61 VGND.n45 9.3005
R5025 VGND.n3235 VGND.n3234 9.3005
R5026 VGND.n3127 VGND.n3126 9.3005
R5027 VGND.n754 VGND.n183 9.3005
R5028 VGND.n729 VGND.n727 9.3005
R5029 VGND.n2568 VGND.n2567 9.3005
R5030 VGND.n1244 VGND.n1218 9.3005
R5031 VGND.n1164 VGND.n7 9.3005
R5032 VGND.n1259 VGND.n1258 9.3005
R5033 VGND.n1263 VGND.n1262 9.3005
R5034 VGND.n1181 VGND.n1180 9.3005
R5035 VGND.t112 VGND.n1397 9.19961
R5036 VGND.n1294 VGND.t97 9.19961
R5037 VGND.t76 VGND.n1381 9.18309
R5038 VGND.t20 VGND.n1278 9.07701
R5039 VGND.n1469 VGND.n1468 8.83211
R5040 VGND.n1212 VGND.n1189 8.73431
R5041 VGND.n1198 VGND.t38 8.63112
R5042 VGND.n1266 VGND.t14 8.63112
R5043 VGND.n1204 VGND.n1203 8.3962
R5044 VGND.n3126 VGND.n167 8.36219
R5045 VGND.n105 VGND.n104 8.33538
R5046 VGND.n3038 VGND.n3037 8.21424
R5047 VGND.n1428 VGND.n1426 8.20035
R5048 VGND.n894 VGND.n893 8.0005
R5049 VGND.t99 VGND.n1287 7.95724
R5050 VGND.n1280 VGND.n1273 7.88469
R5051 VGND.n3118 VGND.n183 7.86418
R5052 VGND.n2567 VGND.n2566 7.74335
R5053 VGND.n1456 VGND.n1390 7.70315
R5054 VGND.n2645 VGND.n766 7.52991
R5055 VGND.n940 VGND.n939 7.52991
R5056 VGND.n756 VGND.n175 7.52991
R5057 VGND.n736 VGND.n185 7.52991
R5058 VGND.n747 VGND.n746 7.52991
R5059 VGND.n773 VGND.n772 7.52991
R5060 VGND.n2625 VGND.n2624 7.52991
R5061 VGND.n192 VGND.n191 7.52991
R5062 VGND.n3132 VGND.n157 7.52991
R5063 VGND.n2851 VGND.n492 7.46717
R5064 VGND.n2296 VGND.n2065 7.46717
R5065 VGND.n2315 VGND.n2314 7.46717
R5066 VGND.n3103 VGND.n3102 7.1223
R5067 VGND.n3102 VGND.n3101 7.1223
R5068 VGND.n3101 VGND.n201 7.1223
R5069 VGND.n204 VGND.n201 7.1223
R5070 VGND.n207 VGND.n204 7.1223
R5071 VGND.n3094 VGND.n207 7.1223
R5072 VGND.n3094 VGND.n3093 7.1223
R5073 VGND.n3093 VGND.n3092 7.1223
R5074 VGND.n3092 VGND.n209 7.1223
R5075 VGND.n215 VGND.n212 7.1223
R5076 VGND.n3085 VGND.n215 7.1223
R5077 VGND.n3085 VGND.n3084 7.1223
R5078 VGND.n3084 VGND.n3083 7.1223
R5079 VGND.n3083 VGND.n217 7.1223
R5080 VGND.n220 VGND.n217 7.1223
R5081 VGND.n223 VGND.n220 7.1223
R5082 VGND.n3077 VGND.n223 7.1223
R5083 VGND.n1439 VGND.n1438 6.83895
R5084 VGND.n3070 VGND.n231 6.72464
R5085 VGND.n231 VGND.n229 6.72464
R5086 VGND.n3068 VGND.n3067 6.72464
R5087 VGND.n3067 VGND.n3066 6.72464
R5088 VGND.n3065 VGND.n3064 6.72464
R5089 VGND.n3066 VGND.n3065 6.72464
R5090 VGND.n238 VGND.n237 6.72464
R5091 VGND.n237 VGND.n236 6.72464
R5092 VGND.n239 VGND.n218 6.72464
R5093 VGND.n236 VGND.n218 6.72464
R5094 VGND.n247 VGND.n246 6.72464
R5095 VGND.n246 VGND.n245 6.72464
R5096 VGND.n244 VGND.n216 6.72464
R5097 VGND.n245 VGND.n244 6.72464
R5098 VGND.n253 VGND.n252 6.72464
R5099 VGND.n254 VGND.n253 6.72464
R5100 VGND.n256 VGND.n255 6.72464
R5101 VGND.n255 VGND.n254 6.72464
R5102 VGND.n264 VGND.n263 6.72464
R5103 VGND.n263 VGND.n262 6.72464
R5104 VGND.n257 VGND.n210 6.72464
R5105 VGND.n262 VGND.n210 6.72464
R5106 VGND.n1100 VGND.n1099 6.72464
R5107 VGND.n1099 VGND.n1098 6.72464
R5108 VGND.n1097 VGND.n208 6.72464
R5109 VGND.n1098 VGND.n1097 6.72464
R5110 VGND.n1109 VGND.n1108 6.72464
R5111 VGND.n1108 VGND.n1107 6.72464
R5112 VGND.n1106 VGND.n1105 6.72464
R5113 VGND.n1107 VGND.n1106 6.72464
R5114 VGND.n1116 VGND.n1115 6.72464
R5115 VGND.n1115 VGND.n1114 6.72464
R5116 VGND.n1117 VGND.n202 6.72464
R5117 VGND.n1114 VGND.n202 6.72464
R5118 VGND.n1127 VGND.n1126 6.72464
R5119 VGND.n1126 VGND.n1125 6.72464
R5120 VGND.n1124 VGND.n200 6.72464
R5121 VGND.n1125 VGND.n1124 6.72464
R5122 VGND.n3076 VGND.n222 6.72464
R5123 VGND.n229 VGND.n222 6.72464
R5124 VGND.n199 VGND.n197 6.72464
R5125 VGND.n1159 VGND.n197 6.72464
R5126 VGND.n1158 VGND.n1157 6.72464
R5127 VGND.n1159 VGND.n1158 6.72464
R5128 VGND.n1534 VGND.n1308 6.6012
R5129 VGND.n1333 VGND.n1308 6.6012
R5130 VGND.n1334 VGND.n1333 6.6012
R5131 VGND.n1523 VGND.n1334 6.6012
R5132 VGND.n1523 VGND.n1522 6.6012
R5133 VGND.n1522 VGND.n1521 6.6012
R5134 VGND.n1521 VGND.n1337 6.6012
R5135 VGND.n1359 VGND.n1337 6.6012
R5136 VGND.n1360 VGND.n1359 6.6012
R5137 VGND.n1510 VGND.n1360 6.6012
R5138 VGND.n1510 VGND.n1509 6.6012
R5139 VGND.n1509 VGND.n1361 6.6012
R5140 VGND.n1499 VGND.n1361 6.6012
R5141 VGND.n1499 VGND.n1498 6.6012
R5142 VGND.n3276 VGND.n10 6.53327
R5143 VGND.n1405 VGND.n1303 6.49846
R5144 VGND.n3236 VGND.n60 6.4522
R5145 VGND.n272 VGND.n271 6.32115
R5146 VGND.n2636 VGND.n2635 6.31912
R5147 VGND.n1194 VGND.n1181 6.1445
R5148 VGND.n1300 VGND.t104 6.13341
R5149 VGND.n1128 VGND.n1091 6.13124
R5150 VGND.n1129 VGND.n1128 6.13124
R5151 VGND.n1129 VGND.n1110 6.13124
R5152 VGND.n1137 VGND.n1110 6.13124
R5153 VGND.n1138 VGND.n1137 6.13124
R5154 VGND.n1139 VGND.n1138 6.13124
R5155 VGND.n1139 VGND.n1093 6.13124
R5156 VGND.n1147 VGND.n1093 6.13124
R5157 VGND.n3045 VGND.n248 6.13124
R5158 VGND.n3053 VGND.n248 6.13124
R5159 VGND.n3054 VGND.n3053 6.13124
R5160 VGND.n3055 VGND.n3054 6.13124
R5161 VGND.n3055 VGND.n232 6.13124
R5162 VGND.n3063 VGND.n232 6.13124
R5163 VGND.n3069 VGND.n3063 6.13124
R5164 VGND.n3071 VGND.n3069 6.13124
R5165 VGND.n1211 VGND.n1190 6.10283
R5166 VGND.n2580 VGND.n958 6.08145
R5167 VGND.n3261 VGND.n3259 6.04885
R5168 VGND.n3110 VGND.n166 5.95912
R5169 VGND.n3134 VGND.n166 5.95912
R5170 VGND.n3134 VGND.n3133 5.95912
R5171 VGND.n3133 VGND.n167 5.95912
R5172 VGND.n3111 VGND.n3110 5.91888
R5173 VGND.n1207 VGND.n1187 5.83948
R5174 VGND.n2627 VGND.n2626 5.83615
R5175 VGND.n2627 VGND.n774 5.83615
R5176 VGND.n2647 VGND.n2646 5.83615
R5177 VGND.n2646 VGND.n762 5.83615
R5178 VGND.n941 VGND.n174 5.83615
R5179 VGND.n3122 VGND.n3121 5.83615
R5180 VGND.n3121 VGND.n176 5.83615
R5181 VGND.n3113 VGND.n176 5.83615
R5182 VGND.n3275 VGND.n11 5.78302
R5183 VGND.n221 VGND.n213 5.77478
R5184 VGND.n1470 VGND.n1469 5.75855
R5185 VGND.n1475 VGND.n1470 5.75855
R5186 VGND.n1476 VGND.n1475 5.75855
R5187 VGND.n1477 VGND.n1476 5.75855
R5188 VGND.n1478 VGND.n1477 5.75855
R5189 VGND.n1479 VGND.n1478 5.75855
R5190 VGND.n1480 VGND.n1479 5.75855
R5191 VGND.n1485 VGND.n1480 5.75855
R5192 VGND.n1486 VGND.n1485 5.75855
R5193 VGND.n1487 VGND.n1486 5.75855
R5194 VGND.n1488 VGND.n1487 5.75855
R5195 VGND.n1492 VGND.n1488 5.75855
R5196 VGND.n1492 VGND.n1491 5.75855
R5197 VGND.n1491 VGND.n13 5.75855
R5198 VGND.n1560 VGND.n1559 5.75855
R5199 VGND.n1559 VGND.n1558 5.75855
R5200 VGND.n1558 VGND.n1283 5.75855
R5201 VGND.n1550 VGND.n1283 5.75855
R5202 VGND.n1550 VGND.n1549 5.75855
R5203 VGND.n1549 VGND.n1548 5.75855
R5204 VGND.n2639 VGND.n731 5.7505
R5205 VGND.n2666 VGND.n731 5.7505
R5206 VGND.n2640 VGND.n732 5.7505
R5207 VGND.n2665 VGND.n732 5.7505
R5208 VGND.n2642 VGND.n733 5.7505
R5209 VGND.n2664 VGND.n733 5.7505
R5210 VGND.n734 VGND.n172 5.7505
R5211 VGND.n2663 VGND.n734 5.7505
R5212 VGND.n735 VGND.n173 5.7505
R5213 VGND.n2662 VGND.n735 5.7505
R5214 VGND.n738 VGND.n737 5.7505
R5215 VGND.n753 VGND.n737 5.7505
R5216 VGND.n751 VGND.n750 5.7505
R5217 VGND.n752 VGND.n751 5.7505
R5218 VGND.n749 VGND.n748 5.7505
R5219 VGND.n748 VGND.n169 5.7505
R5220 VGND.n3131 VGND.n168 5.7505
R5221 VGND.n3131 VGND.n3130 5.7505
R5222 VGND.n830 VGND.n829 5.748
R5223 VGND.n740 VGND.n739 5.748
R5224 VGND.n742 VGND.n741 5.748
R5225 VGND.n1152 VGND.n212 5.6787
R5226 VGND.t88 VGND.n1294 5.65877
R5227 VGND.t51 VGND.n1397 5.65877
R5228 VGND.n2357 VGND.n1014 5.6401
R5229 VGND.n2365 VGND.n2364 5.6401
R5230 VGND.n2373 VGND.n1007 5.6401
R5231 VGND.n2381 VGND.n2380 5.6401
R5232 VGND.n1005 VGND.n1004 5.6401
R5233 VGND.n2389 VGND.n1001 5.6401
R5234 VGND.n1973 VGND.n1081 5.6401
R5235 VGND.n1975 VGND.n1974 5.6401
R5236 VGND.n1982 VGND.n1077 5.6401
R5237 VGND.n1988 VGND.n1074 5.6401
R5238 VGND.n1990 VGND.n1989 5.6401
R5239 VGND.n2000 VGND.n1072 5.6401
R5240 VGND.n1999 VGND.n1070 5.6401
R5241 VGND.n1060 VGND.n1059 5.6401
R5242 VGND.n2325 VGND.n1056 5.6401
R5243 VGND.n2324 VGND.n1057 5.6401
R5244 VGND.n1730 VGND.n1708 5.6401
R5245 VGND.n1726 VGND.n1725 5.6401
R5246 VGND.n1722 VGND.n1721 5.6401
R5247 VGND.n1718 VGND.n1717 5.6401
R5248 VGND.n2951 VGND.n362 5.36011
R5249 VGND.n148 VGND.n123 5.32327
R5250 VGND.n1702 VGND.n1012 5.25991
R5251 VGND.n1246 VGND.n1186 5.23596
R5252 VGND.n2660 VGND.n2659 5.22382
R5253 VGND.n2591 VGND.n2590 5.21817
R5254 VGND.n3274 VGND.n9 5.17867
R5255 VGND.n3045 VGND.n3044 5.17849
R5256 VGND.n1560 VGND.n1281 5.09716
R5257 VGND.n1565 VGND.n1272 5.05856
R5258 VGND.n1564 VGND.n1563 4.99069
R5259 VGND.n1548 VGND.n1297 4.98044
R5260 VGND.n2634 VGND.n2633 4.96999
R5261 VGND.t2 VGND.n1404 4.90692
R5262 VGND.n2358 VGND.n2356 4.87971
R5263 VGND.n1969 VGND.n1968 4.87971
R5264 VGND.n2952 VGND.n359 4.76785
R5265 VGND.n3124 VGND.n3123 4.6505
R5266 VGND.n3277 VGND.n3276 4.6255
R5267 VGND.n1174 VGND.n1 4.54911
R5268 VGND.n2647 VGND.n2644 4.53934
R5269 VGND.n1444 VGND.n1443 4.50187
R5270 VGND.n2677 VGND.n2676 4.5005
R5271 VGND.n3128 VGND.n3127 4.5005
R5272 VGND.n71 VGND.n70 4.5005
R5273 VGND.n75 VGND.n74 4.5005
R5274 VGND.n3193 VGND.n3158 4.5005
R5275 VGND.n3198 VGND.n3197 4.5005
R5276 VGND.n1191 VGND.n1178 4.5005
R5277 VGND.n1244 VGND.n1243 4.5005
R5278 VGND.n67 VGND.n38 4.37945
R5279 VGND.n271 VGND.t108 4.35756
R5280 VGND.n1735 VGND.n1705 4.30941
R5281 VGND.n1155 VGND.n1154 4.26318
R5282 VGND.n1264 VGND.n1263 4.15547
R5283 VGND.n1150 VGND.n268 4.13445
R5284 VGND.n1731 VGND.n1707 4.05595
R5285 VGND.n895 VGND.n894 4.0005
R5286 VGND.n942 VGND.n762 3.98699
R5287 VGND.n1148 VGND.n265 3.9772
R5288 VGND.n3113 VGND.n3112 3.96298
R5289 VGND.t93 VGND.t132 3.92857
R5290 VGND.n3037 VGND.n3036 3.9274
R5291 VGND.n2372 VGND.n2371 3.86585
R5292 VGND.n1981 VGND.n1079 3.86585
R5293 VGND.n1150 VGND.n1149 3.80541
R5294 VGND.n3041 VGND.n268 3.74069
R5295 VGND.n1151 VGND.n267 3.68543
R5296 VGND.n1581 VGND.n970 3.6439
R5297 VGND.n2633 VGND.n779 3.60275
R5298 VGND.n2317 VGND.n1062 3.6005
R5299 VGND.n3043 VGND.n3042 3.53758
R5300 VGND.n2853 VGND.n489 3.52902
R5301 VGND.n2928 VGND.n2927 3.52902
R5302 VGND.n2599 VGND.n947 3.50568
R5303 VGND.n1192 VGND.n1180 3.49908
R5304 VGND.n1967 VGND.n1084 3.49141
R5305 VGND.n3123 VGND.n174 3.48268
R5306 VGND.n133 VGND.n28 3.43465
R5307 VGND.n61 VGND.n48 3.42119
R5308 VGND.t98 VGND.n1404 3.34852
R5309 VGND.n1545 VGND.n1544 3.34148
R5310 VGND.n1230 VGND.t66 3.3065
R5311 VGND.n1230 VGND.t41 3.3065
R5312 VGND.n1221 VGND.t56 3.3065
R5313 VGND.n1221 VGND.t24 3.3065
R5314 VGND.n1222 VGND.t90 3.3065
R5315 VGND.n1222 VGND.t116 3.3065
R5316 VGND.n1224 VGND.t61 3.3065
R5317 VGND.n1224 VGND.t111 3.3065
R5318 VGND.n2678 VGND.n2677 3.30099
R5319 VGND.n145 VGND.n127 3.27855
R5320 VGND.n2672 VGND.n2671 3.22773
R5321 VGND.n1968 VGND.n1083 3.21989
R5322 VGND.n3266 VGND.n19 3.10353
R5323 VGND.n1301 VGND.t58 3.0672
R5324 VGND.n2996 VGND.n2995 3.0005
R5325 VGND.n2955 VGND.n356 2.96248
R5326 VGND.n151 VGND.n150 2.96005
R5327 VGND.n79 VGND.n63 2.88844
R5328 VGND.n3041 VGND.n3040 2.85883
R5329 VGND.n2063 VGND.n1065 2.75742
R5330 VGND.n3234 VGND.n63 2.54637
R5331 VGND.n2671 VGND.n726 2.47089
R5332 VGND.n2713 VGND.n689 2.45829
R5333 VGND.n2744 VGND.n535 2.45829
R5334 VGND.n1462 VGND.n1307 2.4359
R5335 VGND.n424 VGND.n394 2.42922
R5336 VGND.n402 VGND.n400 2.42922
R5337 VGND.n2920 VGND.n2919 2.42922
R5338 VGND.n410 VGND.n408 2.42922
R5339 VGND.n2863 VGND.n2862 2.42922
R5340 VGND.n2859 VGND.n481 2.42922
R5341 VGND.n2858 VGND.n485 2.42922
R5342 VGND.n1852 VGND.n1851 2.42922
R5343 VGND.n1850 VGND.n1849 2.42922
R5344 VGND.n1845 VGND.n1804 2.42922
R5345 VGND.n1844 VGND.n1809 2.42922
R5346 VGND.n1840 VGND.n1839 2.42922
R5347 VGND.n1834 VGND.n1820 2.42922
R5348 VGND.n1830 VGND.n1829 2.42922
R5349 VGND.n1825 VGND.n318 2.42922
R5350 VGND.n2059 VGND.n2058 2.42922
R5351 VGND.n2054 VGND.n1069 2.42922
R5352 VGND.n2053 VGND.n2008 2.42922
R5353 VGND.n2049 VGND.n2048 2.42922
R5354 VGND.n2044 VGND.n2012 2.42922
R5355 VGND.n2039 VGND.n2038 2.42922
R5356 VGND.n2034 VGND.n2021 2.42922
R5357 VGND.n2033 VGND.n2028 2.42922
R5358 VGND.n478 VGND 2.3964
R5359 VGND.n1835 VGND 2.3964
R5360 VGND.n2019 VGND 2.3964
R5361 VGND.n3123 VGND.n3122 2.35397
R5362 VGND.n683 VGND.n680 2.33662
R5363 VGND.n2784 VGND.n2783 2.33662
R5364 VGND.n2673 VGND.n2672 2.3255
R5365 VGND.n952 VGND.n777 2.29818
R5366 VGND.n3039 VGND.n77 2.28623
R5367 VGND.n2316 VGND.n2315 2.28169
R5368 VGND.n1414 VGND.n1407 2.27755
R5369 VGND.n2316 VGND.n1063 2.26512
R5370 VGND.n3125 VGND.n3124 2.2505
R5371 VGND.n3004 VGND.n3003 2.2505
R5372 VGND.n3234 VGND.n3233 2.2505
R5373 VGND.n877 VGND.n874 2.24843
R5374 VGND.n2626 VGND.n779 2.2339
R5375 VGND.n2676 VGND.n721 2.23279
R5376 VGND.n1182 VGND.n1174 2.22861
R5377 VGND.n664 VGND.n663 2.22199
R5378 VGND.n1263 VGND.n1173 2.21202
R5379 VGND.n1751 VGND.n1747 2.19061
R5380 VGND.n1864 VGND.n1858 2.19061
R5381 VGND.n1858 VGND.n1857 2.19061
R5382 VGND.n2246 VGND.n689 2.19061
R5383 VGND.n2725 VGND.n680 2.19061
R5384 VGND.n2744 VGND.n588 2.19061
R5385 VGND.n2783 VGND.n540 2.19061
R5386 VGND.n1935 VGND.n1632 2.19061
R5387 VGND.n2882 VGND.n392 2.19061
R5388 VGND.n2930 VGND.n392 2.19061
R5389 VGND.n3279 VGND.n8 2.18073
R5390 VGND.n2951 VGND.n360 2.15458
R5391 VGND.n1148 VGND.n1147 2.15455
R5392 VGND.n85 VGND.n48 2.15222
R5393 VGND.n2994 VGND.n320 2.14967
R5394 VGND.n1420 VGND.t37 2.14734
R5395 VGND.n1258 VGND.n1173 2.145
R5396 VGND.n1596 VGND.n1595 2.08892
R5397 VGND.n2356 VGND.n1017 2.02027
R5398 VGND.n2679 VGND.n720 2.01471
R5399 VGND.n953 VGND.n360 1.95353
R5400 VGND.n1897 VGND.n1655 1.93989
R5401 VGND.n1697 VGND.n1696 1.93989
R5402 VGND.n1661 VGND.n1657 1.93989
R5403 VGND.n1690 VGND.n1662 1.93989
R5404 VGND.n1689 VGND.n1663 1.93989
R5405 VGND.n1683 VGND.n1682 1.93989
R5406 VGND.n1668 VGND.n1665 1.93989
R5407 VGND.n1676 VGND.n1669 1.93989
R5408 VGND.n1675 VGND.n1671 1.93989
R5409 VGND.n1637 VGND.n1636 1.93989
R5410 VGND.n1926 VGND.n1638 1.93989
R5411 VGND.n1925 VGND.n1923 1.93989
R5412 VGND.n1922 VGND.n1639 1.93989
R5413 VGND.n1919 VGND.n1918 1.93989
R5414 VGND.n1742 VGND.n1640 1.93989
R5415 VGND.n1912 VGND.n1648 1.93989
R5416 VGND.n1911 VGND.n1649 1.93989
R5417 VGND.n1908 VGND.n1907 1.93989
R5418 VGND.n1961 VGND.n1603 1.93989
R5419 VGND.n1960 VGND.n1604 1.93989
R5420 VGND.n1956 VGND.n1955 1.93989
R5421 VGND.n1611 VGND.n1607 1.93989
R5422 VGND.n1949 VGND.n1612 1.93989
R5423 VGND.n1948 VGND.n1613 1.93989
R5424 VGND.n1944 VGND.n1943 1.93989
R5425 VGND.n1620 VGND.n1617 1.93989
R5426 VGND.n1937 VGND.n1626 1.93989
R5427 VGND.n3236 VGND.n3235 1.93153
R5428 VGND.n686 VGND.n683 1.92293
R5429 VGND.n2785 VGND.n2784 1.92293
R5430 VGND.n2713 VGND.n686 1.8986
R5431 VGND.n2785 VGND.n535 1.8986
R5432 VGND.n2635 VGND.n2634 1.85779
R5433 VGND.n2989 VGND.n2988 1.85174
R5434 VGND.n336 VGND.n331 1.85174
R5435 VGND.n2972 VGND.n334 1.85174
R5436 VGND.n2966 VGND.n2965 1.85174
R5437 VGND.n2355 VGND.n1022 1.84993
R5438 VGND.n942 VGND.n941 1.84966
R5439 VGND.n1193 VGND.n1192 1.84749
R5440 VGND.n2589 VGND.n2588 1.84721
R5441 VGND.n1541 VGND.n1304 1.83816
R5442 VGND.n3232 VGND.n3231 1.81528
R5443 VGND.n3287 VGND.n1 1.80047
R5444 VGND.n3284 VGND.n4 1.79699
R5445 VGND.n1214 VGND.n1213 1.79521
R5446 VGND.n3219 VGND.n3218 1.77828
R5447 VGND.n2374 VGND.n2372 1.77476
R5448 VGND.n341 VGND.n339 1.7724
R5449 VGND.n3026 VGND.n3025 1.7505
R5450 VGND.n3020 VGND.n290 1.7505
R5451 VGND.n811 VGND.n291 1.7505
R5452 VGND.n825 VGND.n823 1.7505
R5453 VGND.n308 VGND.n306 1.7505
R5454 VGND.n3009 VGND.n310 1.7505
R5455 VGND.n3258 VGND.n26 1.74306
R5456 VGND.n1250 VGND.n1177 1.73997
R5457 VGND.n2683 VGND.n2682 1.73791
R5458 VGND.n976 VGND.n972 1.7358
R5459 VGND.n2589 VGND.n730 1.73158
R5460 VGND.n1751 VGND.n1700 1.70392
R5461 VGND.n1888 VGND.n1887 1.70392
R5462 VGND.n1884 VGND.n1762 1.70392
R5463 VGND.n1767 VGND.n1763 1.70392
R5464 VGND.n1878 VGND.n1774 1.70392
R5465 VGND.n1874 VGND.n1873 1.70392
R5466 VGND.n1870 VGND.n1782 1.70392
R5467 VGND.n2180 VGND.n692 1.70392
R5468 VGND.n2707 VGND.n695 1.70392
R5469 VGND.n2199 VGND.n2181 1.70392
R5470 VGND.n2207 VGND.n2185 1.70392
R5471 VGND.n2196 VGND.n2189 1.70392
R5472 VGND.n2193 VGND.n982 1.70392
R5473 VGND.n2428 VGND.n2426 1.70392
R5474 VGND.n2295 VGND.n2069 1.70392
R5475 VGND.n2292 VGND.n2075 1.70392
R5476 VGND.n2288 VGND.n2287 1.70392
R5477 VGND.n2284 VGND.n2080 1.70392
R5478 VGND.n2108 VGND.n2081 1.70392
R5479 VGND.n2277 VGND.n2115 1.70392
R5480 VGND.n2273 VGND.n2272 1.70392
R5481 VGND.n2269 VGND.n2126 1.70392
R5482 VGND.n2247 VGND.n2127 1.70392
R5483 VGND.n2850 VGND.n495 1.70392
R5484 VGND.n2846 VGND.n2845 1.70392
R5485 VGND.n2841 VGND.n503 1.70392
R5486 VGND.n506 VGND.n504 1.70392
R5487 VGND.n2811 VGND.n512 1.70392
R5488 VGND.n2805 VGND.n2804 1.70392
R5489 VGND.n2800 VGND.n521 1.70392
R5490 VGND.n524 VGND.n522 1.70392
R5491 VGND.n2792 VGND.n529 1.70392
R5492 VGND.n2771 VGND.n568 1.70392
R5493 VGND.n2768 VGND.n2767 1.70392
R5494 VGND.n2752 VGND.n576 1.70392
R5495 VGND.n2762 VGND.n578 1.70392
R5496 VGND.n2757 VGND.n580 1.70392
R5497 VGND.n2473 VGND.n2472 1.70392
R5498 VGND.n2477 VGND.n2476 1.70392
R5499 VGND.n1632 VGND.n432 1.70392
R5500 VGND.n2908 VGND.n2907 1.70392
R5501 VGND.n450 VGND.n442 1.70392
R5502 VGND.n2902 VGND.n447 1.70392
R5503 VGND.n449 VGND.n448 1.70392
R5504 VGND.n2897 VGND.n457 1.70392
R5505 VGND.n2890 VGND.n2889 1.70392
R5506 VGND.n1252 VGND.n1251 1.69667
R5507 VGND.n1409 VGND.n1407 1.69277
R5508 VGND.n3203 VGND.n3153 1.68289
R5509 VGND.n954 VGND.n953 1.68066
R5510 VGND.n2984 VGND.n327 1.66662
R5511 VGND.n2983 VGND.n328 1.66662
R5512 VGND.n2950 VGND.n367 1.66662
R5513 VGND.t130 VGND.n1301 1.66381
R5514 VGND.n1413 VGND.n9 1.66095
R5515 VGND.n2699 VGND.n2698 1.6499
R5516 VGND.n741 VGND.n740 1.648
R5517 VGND.n1248 VGND.n1181 1.62685
R5518 VGND.n3280 VGND.n7 1.61213
R5519 VGND.n2869 VGND.n2868 1.60871
R5520 VGND.n1246 VGND.n1245 1.59631
R5521 VGND.t52 VGND.n299 1.58922
R5522 VGND.n1581 VGND.t109 1.58479
R5523 VGND.n1707 VGND.n1706 1.58466
R5524 VGND.n1670 VGND.n282 1.5755
R5525 VGND.n1563 VGND.n1274 1.57523
R5526 VGND.n1555 VGND.n1274 1.57523
R5527 VGND.n1555 VGND.n1554 1.57523
R5528 VGND.n1554 VGND.n1553 1.57523
R5529 VGND.n1545 VGND.n1302 1.57523
R5530 VGND.n1422 VGND.n1420 1.55836
R5531 VGND.n1898 VGND.n1897 1.55202
R5532 VGND.n1697 VGND.n1655 1.55202
R5533 VGND.n1696 VGND.n1657 1.55202
R5534 VGND.n1662 VGND.n1661 1.55202
R5535 VGND.n1690 VGND.n1689 1.55202
R5536 VGND.n1683 VGND.n1663 1.55202
R5537 VGND.n1682 VGND.n1665 1.55202
R5538 VGND.n1669 VGND.n1668 1.55202
R5539 VGND.n1676 VGND.n1675 1.55202
R5540 VGND.n1636 VGND.n1627 1.55202
R5541 VGND.n1638 VGND.n1637 1.55202
R5542 VGND.n1926 VGND.n1925 1.55202
R5543 VGND.n1923 VGND.n1922 1.55202
R5544 VGND.n1919 VGND.n1639 1.55202
R5545 VGND.n1918 VGND.n1640 1.55202
R5546 VGND.n1912 VGND.n1911 1.55202
R5547 VGND.n1908 VGND.n1649 1.55202
R5548 VGND.n1603 VGND.n1084 1.55202
R5549 VGND.n1961 VGND.n1960 1.55202
R5550 VGND.n1956 VGND.n1604 1.55202
R5551 VGND.n1955 VGND.n1607 1.55202
R5552 VGND.n1612 VGND.n1611 1.55202
R5553 VGND.n1949 VGND.n1948 1.55202
R5554 VGND.n1944 VGND.n1613 1.55202
R5555 VGND.n1943 VGND.n1617 1.55202
R5556 VGND.n1626 VGND.n1620 1.55202
R5557 VGND.n1574 VGND.n1573 1.54681
R5558 VGND.n2445 VGND.n972 1.54681
R5559 VGND.n2698 VGND.n705 1.54681
R5560 VGND.n2592 VGND.n2586 1.54488
R5561 VGND.n3251 VGND.n33 1.53643
R5562 VGND.n3251 VGND.n3250 1.53557
R5563 VGND.n1747 VGND.n1650 1.53358
R5564 VGND.n1936 VGND.n1935 1.53358
R5565 VGND.n1738 VGND.n1075 1.52129
R5566 VGND.n2315 VGND.n1060 1.52129
R5567 VGND.n743 VGND.n274 1.50813
R5568 VGND.n3252 VGND.n32 1.48623
R5569 VGND.n74 VGND.n73 1.48012
R5570 VGND.n1125 VGND.n1122 1.45636
R5571 VGND.n1114 VGND.n1112 1.45636
R5572 VGND.n1107 VGND.n1103 1.45636
R5573 VGND.n1098 VGND.n1095 1.45636
R5574 VGND.n262 VGND.n260 1.45636
R5575 VGND.n254 VGND.n250 1.45636
R5576 VGND.n245 VGND.n242 1.45636
R5577 VGND.n3066 VGND.n228 1.45636
R5578 VGND.n3280 VGND.n3279 1.45587
R5579 VGND.n1594 VGND.n1585 1.45523
R5580 VGND.n115 VGND.n34 1.45347
R5581 VGND.n1152 VGND.n209 1.44411
R5582 VGND.n236 VGND.n234 1.44145
R5583 VGND.n1570 VGND.n1002 1.42654
R5584 VGND.n3015 VGND.n3014 1.4255
R5585 VGND.n1757 VGND.n1746 1.41191
R5586 VGND.n2677 VGND.n722 1.40335
R5587 VGND.n68 VGND.n66 1.40196
R5588 VGND.n1205 VGND.n1193 1.36456
R5589 VGND.n1743 VGND.n1648 1.35808
R5590 VGND.n1259 VGND.n1175 1.35794
R5591 VGND.n2699 VGND.n704 1.35782
R5592 VGND.n835 VGND.n812 1.3505
R5593 VGND.n1591 VGND.n1590 1.34787
R5594 VGND.n976 VGND.n704 1.34063
R5595 VGND.n1735 VGND.n1734 1.33119
R5596 VGND.n1302 VGND.n1290 1.33051
R5597 VGND.n3255 VGND.n3254 1.32811
R5598 VGND.n3178 VGND.n3173 1.3278
R5599 VGND.n3164 VGND.n3163 1.3278
R5600 VGND.n2989 VGND.n323 1.32281
R5601 VGND.n878 VGND.n877 1.32281
R5602 VGND.n3178 VGND.n80 1.31506
R5603 VGND.n3163 VGND.n3150 1.31505
R5604 VGND.n3216 VGND.n45 1.31382
R5605 VGND.n3198 VGND.n3158 1.31136
R5606 VGND.n3282 VGND.n6 1.30959
R5607 VGND.n2644 VGND.n774 1.29731
R5608 VGND.n1621 VGND.n434 1.29023
R5609 VGND.n1542 VGND.n1541 1.27937
R5610 VGND.n3130 VGND.n3129 1.27722
R5611 VGND.n2594 VGND.n951 1.27684
R5612 VGND.n285 VGND.n282 1.2755
R5613 VGND.n3004 VGND.n311 1.2755
R5614 VGND.n1573 VGND.n998 1.27191
R5615 VGND.n2396 VGND.n2395 1.27191
R5616 VGND.n999 VGND.n994 1.27191
R5617 VGND.n2404 VGND.n2402 1.27191
R5618 VGND.n2403 VGND.n992 1.27191
R5619 VGND.n991 VGND.n987 1.27191
R5620 VGND.n2419 VGND.n2417 1.27191
R5621 VGND.n2418 VGND.n971 1.27191
R5622 VGND.n710 VGND.n705 1.27191
R5623 VGND.n2692 VGND.n2691 1.27191
R5624 VGND.n2687 VGND.n711 1.27191
R5625 VGND.n2388 VGND.n1002 1.26783
R5626 VGND.n2064 VGND.n1064 1.26783
R5627 VGND.n2356 VGND.n1016 1.26783
R5628 VGND VGND.n2410 1.25473
R5629 VGND.n3228 VGND.n44 1.2487
R5630 VGND.n1210 VGND.n1206 1.24255
R5631 VGND.n37 VGND.n33 1.22178
R5632 VGND.n3250 VGND.n3249 1.22178
R5633 VGND.n3253 VGND.n31 1.21824
R5634 VGND.n2853 VGND.n2852 1.21723
R5635 VGND.n2927 VGND.n397 1.21723
R5636 VGND.n68 VGND.n67 1.2151
R5637 VGND.n3273 VGND.n12 1.21186
R5638 VGND.n1538 VGND.n1537 1.2035
R5639 VGND.n2595 VGND.n2594 1.17858
R5640 VGND.n2595 VGND.n726 1.17858
R5641 VGND.n3129 VGND.n3128 1.17339
R5642 VGND.n3038 VGND.n274 1.16698
R5643 VGND.n69 VGND.n68 1.163
R5644 VGND.n3172 VGND.n3171 1.163
R5645 VGND.n3203 VGND.n3202 1.163
R5646 VGND.n3208 VGND.n3207 1.163
R5647 VGND.n3226 VGND.n3225 1.163
R5648 VGND.n3218 VGND.n3217 1.163
R5649 VGND.n3184 VGND.n3183 1.163
R5650 VGND.n3191 VGND.n3190 1.163
R5651 VGND.n2686 VGND.n714 1.16178
R5652 VGND.n1208 VGND.n1207 1.15586
R5653 VGND.n41 VGND.n40 1.13312
R5654 VGND.n72 VGND.n64 1.1305
R5655 VGND.n1232 VGND.n1231 1.12069
R5656 VGND.n1787 VGND.n1783 1.11989
R5657 VGND.n2878 VGND.n2872 1.11989
R5658 VGND.n2552 VGND.n2455 1.11787
R5659 VGND.n3194 VGND.n3193 1.10831
R5660 VGND.n3160 VGND.n3159 1.10831
R5661 VGND.n3181 VGND.n3180 1.10831
R5662 VGND.n2669 VGND.n727 1.10572
R5663 VGND.n2565 VGND.n2564 1.09556
R5664 VGND.n1540 VGND.n1539 1.09525
R5665 VGND.n3195 VGND.n3152 1.0952
R5666 VGND.n3230 VGND.n77 1.0951
R5667 VGND.n3174 VGND.n78 1.09141
R5668 VGND.n3205 VGND.n3151 1.0914
R5669 VGND.n1253 VGND.n1252 1.08952
R5670 VGND.n723 VGND.n722 1.08232
R5671 VGND.n1229 VGND.n1228 1.08223
R5672 VGND.n3140 VGND.n156 1.07163
R5673 VGND.n1249 VGND.n1179 1.063
R5674 VGND.n2483 VGND.n2459 1.06256
R5675 VGND.n323 VGND.n320 1.05835
R5676 VGND.n878 VGND.n345 1.05835
R5677 VGND.n1233 VGND.n1229 1.05338
R5678 VGND.n978 VGND.n969 1.04689
R5679 VGND.n122 VGND.n121 1.03492
R5680 VGND.n3259 VGND.n3258 1.03383
R5681 VGND.n123 VGND.n122 1.03383
R5682 VGND.n3039 VGND.n3038 1.0281
R5683 VGND.n1227 VGND.n1226 1.02454
R5684 VGND.n3127 VGND.n170 1.02174
R5685 VGND.n1228 VGND.n1227 1.01733
R5686 VGND.n1593 VGND.n1588 0.999039
R5687 VGND.n2559 VGND.n2455 0.996178
R5688 VGND.n2486 VGND.n2483 0.996178
R5689 VGND.n1408 VGND.n1304 0.994585
R5690 VGND.n1305 VGND.n1290 0.983286
R5691 VGND.n2977 VGND.n2976 0.979012
R5692 VGND.n1411 VGND.n1410 0.978812
R5693 VGND.n3026 VGND.n285 0.9755
R5694 VGND.n796 VGND.n288 0.9755
R5695 VGND.n3008 VGND.n311 0.9755
R5696 VGND.n2351 VGND.n2350 0.973884
R5697 VGND.n1030 VGND.n1027 0.973884
R5698 VGND.n2345 VGND.n1032 0.973884
R5699 VGND.n2341 VGND.n2340 0.973884
R5700 VGND.n2333 VGND.n1038 0.973884
R5701 VGND.n2232 VGND.n2231 0.973884
R5702 VGND.n2239 VGND.n2238 0.973884
R5703 VGND.n2251 VGND.n2215 0.973884
R5704 VGND.n2725 VGND.n681 0.973884
R5705 VGND.n2262 VGND.n2261 0.973884
R5706 VGND.n2152 VGND.n2151 0.973884
R5707 VGND.n2170 VGND.n2139 0.973884
R5708 VGND.n2732 VGND.n2731 0.973884
R5709 VGND.n2737 VGND.n2736 0.973884
R5710 VGND.n2158 VGND.n592 0.973884
R5711 VGND.n546 VGND.n540 0.973884
R5712 VGND.n2778 VGND.n2777 0.973884
R5713 VGND.n631 VGND.n630 0.973884
R5714 VGND.n637 VGND.n636 0.973884
R5715 VGND.n621 VGND.n615 0.973884
R5716 VGND.n654 VGND.n612 0.973884
R5717 VGND.n657 VGND.n610 0.973884
R5718 VGND.n659 VGND.n349 0.973884
R5719 VGND.n370 VGND.n361 0.967441
R5720 VGND.n1225 VGND.n1216 0.964541
R5721 VGND.t7 VGND.n221 0.961828
R5722 VGND.n3044 VGND.n265 0.953251
R5723 VGND.n2227 VGND 0.949549
R5724 VGND VGND.n2143 0.949549
R5725 VGND VGND.n619 0.949549
R5726 VGND.n3208 VGND.n82 0.948648
R5727 VGND.n2668 VGND.n2667 0.932326
R5728 VGND.n2634 VGND.n775 0.931491
R5729 VGND.n2512 VGND.n2504 0.923023
R5730 VGND.n2510 VGND.n2509 0.923023
R5731 VGND.n3246 VGND.n3245 0.922756
R5732 VGND.n3257 VGND.n19 0.910217
R5733 VGND.n3242 VGND.n45 0.910039
R5734 VGND.n3040 VGND.n273 0.905089
R5735 VGND.n664 VGND.n356 0.899674
R5736 VGND.n3288 VGND.n3287 0.89249
R5737 VGND.n3258 VGND.n3257 0.884429
R5738 VGND.n2296 VGND.n397 0.876546
R5739 VGND.n2852 VGND.n2851 0.876546
R5740 VGND.n2551 VGND.n2459 0.874484
R5741 VGND.n2978 VGND.n2977 0.873227
R5742 VGND.n1592 VGND.n722 0.868655
R5743 VGND.n3243 VGND.n44 0.864562
R5744 VGND.n2552 VGND.n2551 0.863421
R5745 VGND.n2660 VGND.n183 0.861487
R5746 VGND.n122 VGND.n27 0.858936
R5747 VGND.n102 VGND.n97 0.850998
R5748 VGND.n831 VGND.n830 0.8505
R5749 VGND.n3256 VGND.n28 0.849283
R5750 VGND.n127 VGND.n27 0.847459
R5751 VGND.n2818 VGND.n2817 0.846781
R5752 VGND.n739 VGND.n358 0.84349
R5753 VGND.n2350 VGND.n2349 0.827876
R5754 VGND.n2346 VGND.n1030 0.827876
R5755 VGND.n1034 VGND.n1032 0.827876
R5756 VGND.n2340 VGND.n1036 0.827876
R5757 VGND.n2333 VGND.n2332 0.827876
R5758 VGND.n2227 VGND.n2220 0.827876
R5759 VGND.n2231 VGND.n2219 0.827876
R5760 VGND.n2238 VGND.n2237 0.827876
R5761 VGND.n2251 VGND.n2250 0.827876
R5762 VGND.n2263 VGND.n681 0.827876
R5763 VGND.n2261 VGND.n2131 0.827876
R5764 VGND.n2153 VGND.n2152 0.827876
R5765 VGND.n2170 VGND.n2169 0.827876
R5766 VGND.n2175 VGND.n2138 0.827876
R5767 VGND.n2143 VGND.n602 0.827876
R5768 VGND.n2732 VGND.n594 0.827876
R5769 VGND.n2736 VGND.n596 0.827876
R5770 VGND.n2159 VGND.n2158 0.827876
R5771 VGND.n546 VGND.n543 0.827876
R5772 VGND.n2777 VGND.n545 0.827876
R5773 VGND.n630 VGND.n629 0.827876
R5774 VGND.n636 VGND.n634 0.827876
R5775 VGND.n647 VGND.n615 0.827876
R5776 VGND.n619 VGND.n613 0.827876
R5777 VGND.n654 VGND.n653 0.827876
R5778 VGND.n658 VGND.n657 0.827876
R5779 VGND.n2961 VGND.n349 0.827876
R5780 VGND.n2869 VGND.n469 0.821013
R5781 VGND.n2577 VGND.n2576 0.819169
R5782 VGND.n2453 VGND.n964 0.819169
R5783 VGND.n2560 VGND.n2454 0.819169
R5784 VGND.n2487 VGND.n2486 0.819169
R5785 VGND.n2540 VGND.n2539 0.819169
R5786 VGND.n2536 VGND.n2535 0.819169
R5787 VGND.n2532 VGND.n2488 0.819169
R5788 VGND.n2531 VGND.n2489 0.819169
R5789 VGND.n2525 VGND.n2524 0.819169
R5790 VGND.n2522 VGND.n2521 0.819169
R5791 VGND.n2520 VGND.n2517 0.819169
R5792 VGND.n2951 VGND.n361 0.814262
R5793 VGND.n2498 VGND 0.808106
R5794 VGND.n2597 VGND.n2596 0.797287
R5795 VGND.n2952 VGND.n2951 0.784173
R5796 VGND.n796 VGND.n286 0.7755
R5797 VGND.n2951 VGND.n2950 0.767442
R5798 VGND.n3200 VGND.n3199 0.763261
R5799 VGND.n1210 VGND.n1209 0.761584
R5800 VGND.n2667 VGND.n2666 0.756589
R5801 VGND.n2255 VGND.n2179 0.754873
R5802 VGND.n566 VGND.n534 0.754873
R5803 VGND.n3128 VGND.n3125 0.753367
R5804 VGND.n3184 VGND.n3166 0.747945
R5805 VGND.n1409 VGND.n1305 0.727693
R5806 VGND.n77 VGND.n8 0.718542
R5807 VGND.n3036 VGND.n275 0.716113
R5808 VGND.n2818 VGND.n342 0.71455
R5809 VGND.n663 VGND.n367 0.71455
R5810 VGND.n3202 VGND.n3149 0.711611
R5811 VGND VGND.n3039 0.710753
R5812 VGND.n3281 VGND.n3 0.710675
R5813 VGND.n125 VGND.n29 0.702939
R5814 VGND.n73 VGND.n70 0.69887
R5815 VGND.n743 VGND.n742 0.682643
R5816 VGND.n968 VGND.n967 0.675349
R5817 VGND.n2179 VGND.n686 0.657534
R5818 VGND.n979 VGND.n969 0.657534
R5819 VGND.n2785 VGND.n534 0.657534
R5820 VGND.n1253 VGND.n2 0.653124
R5821 VGND.n1400 VGND.n1303 0.649544
R5822 VGND.n72 VGND.n71 0.643
R5823 VGND.n1215 VGND.n1187 0.638661
R5824 VGND.t107 VGND.n299 0.636287
R5825 VGND.n2995 VGND.n2994 0.6255
R5826 VGND.n2565 VGND.n2450 0.608865
R5827 VGND.n2176 VGND.n2175 0.608865
R5828 VGND.n2956 VGND.n355 0.608764
R5829 VGND.n3162 VGND.n3147 0.607397
R5830 VGND.n1078 VGND.n1063 0.591269
R5831 VGND.n1787 VGND.n468 0.589305
R5832 VGND.n2872 VGND.n2871 0.589305
R5833 VGND.n1790 VGND.n1787 0.58453
R5834 VGND.n2296 VGND.n2295 0.58453
R5835 VGND.n2851 VGND.n2850 0.58453
R5836 VGND.n2885 VGND.n2872 0.58453
R5837 VGND.n2679 VGND.n2678 0.58246
R5838 VGND.n3251 VGND.n34 0.58175
R5839 VGND.n3248 VGND.n38 0.58175
R5840 VGND.n1245 VGND.n1216 0.578692
R5841 VGND.n3278 VGND.n3277 0.577096
R5842 VGND.n3217 VGND.n76 0.563
R5843 VGND.n69 VGND.n42 0.563
R5844 VGND.n3192 VGND.n3191 0.563
R5845 VGND.n3204 VGND.n3203 0.563
R5846 VGND.n3190 VGND.n3188 0.561084
R5847 VGND.n1857 VGND.n1856 0.560196
R5848 VGND.n2930 VGND.n2929 0.560196
R5849 VGND.n1544 VGND.n1543 0.548389
R5850 VGND.n2448 VGND.n969 0.544527
R5851 VGND.n3182 VGND.n3181 0.542167
R5852 VGND.n3182 VGND.n3159 0.540273
R5853 VGND.n105 VGND.n38 0.539447
R5854 VGND.n2667 VGND.n730 0.536723
R5855 VGND.n2449 VGND.n776 0.535881
R5856 VGND.n1411 VGND.n1407 0.534082
R5857 VGND.n2988 VGND.n324 0.529426
R5858 VGND.n2984 VGND.n2983 0.529426
R5859 VGND.n331 VGND.n330 0.529426
R5860 VGND.n2976 VGND.n334 0.529426
R5861 VGND.n2972 VGND.n2971 0.529426
R5862 VGND.n342 VGND.n341 0.529426
R5863 VGND.n2966 VGND.n344 0.529426
R5864 VGND.n2965 VGND.n345 0.529426
R5865 VGND.n1583 VGND.n1582 0.526527
R5866 VGND.n424 VGND.n400 0.525628
R5867 VGND.n2920 VGND.n402 0.525628
R5868 VGND.n2919 VGND.n408 0.525628
R5869 VGND.n469 VGND.n410 0.525628
R5870 VGND.n2863 VGND.n478 0.525628
R5871 VGND.n2862 VGND.n481 0.525628
R5872 VGND.n2859 VGND.n2858 0.525628
R5873 VGND.n487 VGND.n485 0.525628
R5874 VGND.n1851 VGND.n1850 0.525628
R5875 VGND.n1849 VGND.n1804 0.525628
R5876 VGND.n1845 VGND.n1844 0.525628
R5877 VGND.n1840 VGND.n1809 0.525628
R5878 VGND.n1835 VGND.n1834 0.525628
R5879 VGND.n1830 VGND.n1820 0.525628
R5880 VGND.n1829 VGND.n1825 0.525628
R5881 VGND.n2997 VGND.n318 0.525628
R5882 VGND.n2058 VGND.n1069 0.525628
R5883 VGND.n2054 VGND.n2053 0.525628
R5884 VGND.n2049 VGND.n2008 0.525628
R5885 VGND.n2048 VGND.n2012 0.525628
R5886 VGND.n2039 VGND.n2019 0.525628
R5887 VGND.n2038 VGND.n2021 0.525628
R5888 VGND.n2034 VGND.n2033 0.525628
R5889 VGND.n2028 VGND.n395 0.525628
R5890 VGND.n1670 VGND.n276 0.5255
R5891 VGND.n3244 VGND.n43 0.525121
R5892 VGND.n3181 VGND.n43 0.525121
R5893 VGND.n2511 VGND.n2506 0.522949
R5894 VGND.n2587 VGND.n775 0.519538
R5895 VGND.n1746 VGND.n1745 0.517167
R5896 VGND.n2566 VGND.n2565 0.517167
R5897 VGND.n1741 VGND.n434 0.517167
R5898 VGND.n1900 VGND.n1650 0.511527
R5899 VGND.n1936 VGND.n1628 0.511527
R5900 VGND.n3192 VGND.n3159 0.50997
R5901 VGND.n3193 VGND.n3192 0.508076
R5902 VGND.n2513 VGND.n2502 0.504934
R5903 VGND.n1968 VGND.n1967 0.504742
R5904 VGND.n71 VGND.n42 0.504288
R5905 VGND.n3244 VGND.n42 0.502394
R5906 VGND.n3025 VGND.n286 0.5005
R5907 VGND.n290 VGND.n288 0.5005
R5908 VGND.n812 VGND.n811 0.5005
R5909 VGND.n828 VGND.n823 0.5005
R5910 VGND.n825 VGND.n305 0.5005
R5911 VGND.n3014 VGND.n306 0.5005
R5912 VGND.n3009 VGND.n3008 0.5005
R5913 VGND.n3172 VGND.n43 0.5005
R5914 VGND.n3227 VGND.n3226 0.5005
R5915 VGND.n3207 VGND.n3206 0.5005
R5916 VGND.n3183 VGND.n3182 0.5005
R5917 VGND.n2596 VGND.n2595 0.489974
R5918 VGND.n2436 VGND.n704 0.487192
R5919 VGND.n2717 VGND.n686 0.487192
R5920 VGND.n2786 VGND.n2785 0.487192
R5921 VGND.n2551 VGND.n2550 0.487192
R5922 VGND.n3285 VGND.n3 0.486062
R5923 VGND.n3206 VGND.n78 0.477785
R5924 VGND.n3206 VGND.n3205 0.477153
R5925 VGND.n3227 VGND.n78 0.46449
R5926 VGND.n3228 VGND.n3227 0.464045
R5927 VGND.n1543 VGND.n1542 0.463665
R5928 VGND.n1893 VGND.n1700 0.462857
R5929 VGND.n1758 VGND.n1757 0.462857
R5930 VGND.n1887 VGND.n1761 0.462857
R5931 VGND.n1884 VGND.n1883 0.462857
R5932 VGND.n1879 VGND.n1767 0.462857
R5933 VGND.n1778 VGND.n1774 0.462857
R5934 VGND.n1873 VGND.n1781 0.462857
R5935 VGND.n1870 VGND.n1869 0.462857
R5936 VGND.n1865 VGND.n1790 0.462857
R5937 VGND.n2256 VGND.n2255 0.462857
R5938 VGND.n2180 VGND.n694 0.462857
R5939 VGND.n2200 VGND.n695 0.462857
R5940 VGND.n2197 VGND.n2181 0.462857
R5941 VGND.n2207 VGND.n2206 0.462857
R5942 VGND.n2190 VGND.n2189 0.462857
R5943 VGND.n2429 VGND.n982 0.462857
R5944 VGND.n2426 VGND.n980 0.462857
R5945 VGND.n2435 VGND.n978 0.462857
R5946 VGND.n2072 VGND.n2069 0.462857
R5947 VGND.n2077 VGND.n2075 0.462857
R5948 VGND.n2287 VGND.n2079 0.462857
R5949 VGND.n2278 VGND.n2108 0.462857
R5950 VGND.n2120 VGND.n2115 0.462857
R5951 VGND.n2272 VGND.n2123 0.462857
R5952 VGND.n2269 VGND.n2268 0.462857
R5953 VGND.n2247 VGND.n685 0.462857
R5954 VGND.n497 VGND.n495 0.462857
R5955 VGND.n2845 VGND.n500 0.462857
R5956 VGND.n2841 VGND.n2840 0.462857
R5957 VGND.n514 VGND.n512 0.462857
R5958 VGND.n2804 VGND.n517 0.462857
R5959 VGND.n2800 VGND.n2799 0.462857
R5960 VGND.n2793 VGND.n524 0.462857
R5961 VGND.n531 VGND.n529 0.462857
R5962 VGND.n2772 VGND.n566 0.462857
R5963 VGND.n571 VGND.n568 0.462857
R5964 VGND.n2767 VGND.n574 0.462857
R5965 VGND.n2758 VGND.n576 0.462857
R5966 VGND.n2762 VGND.n2761 0.462857
R5967 VGND.n2470 VGND.n580 0.462857
R5968 VGND.n2473 VGND.n2462 0.462857
R5969 VGND.n2476 VGND.n2466 0.462857
R5970 VGND.n2564 VGND.n2451 0.462857
R5971 VGND.n2913 VGND.n432 0.462857
R5972 VGND.n1621 VGND.n437 0.462857
R5973 VGND.n2907 VGND.n440 0.462857
R5974 VGND.n446 VGND.n442 0.462857
R5975 VGND.n2902 VGND.n2901 0.462857
R5976 VGND.n2898 VGND.n449 0.462857
R5977 VGND.n459 VGND.n457 0.462857
R5978 VGND.n2889 VGND.n463 0.462857
R5979 VGND.n2885 VGND.n2884 0.462857
R5980 VGND.n3229 VGND.n76 0.461026
R5981 VGND.n2500 VGND.n370 0.460036
R5982 VGND.n2316 VGND.n2064 0.459987
R5983 VGND.n121 VGND.n120 0.452423
R5984 VGND.n1741 VGND.n1740 0.451467
R5985 VGND.n3205 VGND.n3204 0.450893
R5986 VGND.n2638 VGND.n775 0.448409
R5987 VGND.n2594 VGND.n2593 0.447421
R5988 VGND.n3204 VGND.n3152 0.445463
R5989 VGND.n1594 VGND.n1593 0.44374
R5990 VGND.n1017 VGND.n1009 0.438523
R5991 VGND.n2590 VGND.n950 0.437448
R5992 VGND.n1165 VGND.n1164 0.436864
R5993 VGND.n2566 VGND.n2449 0.433025
R5994 VGND.n2568 VGND.n963 0.431961
R5995 VGND.n26 VGND.n25 0.428385
R5996 VGND.n2064 VGND.n2063 0.427167
R5997 VGND.n3217 VGND.n3216 0.426133
R5998 VGND.n1175 VGND.n2 0.425272
R5999 VGND.n3257 VGND.n3256 0.424111
R6000 VGND.n3286 VGND.n3285 0.423372
R6001 VGND.n70 VGND.n37 0.4221
R6002 VGND.n3183 VGND.n3173 0.422012
R6003 VGND.n3183 VGND.n3164 0.420558
R6004 VGND.n3242 VGND.n36 0.418263
R6005 VGND.n3256 VGND.n27 0.417167
R6006 VGND.n1745 VGND.n275 0.414879
R6007 VGND.n2912 VGND.n434 0.414188
R6008 VGND.n1736 VGND.n1704 0.410297
R6009 VGND.n3172 VGND.n36 0.40893
R6010 VGND.n3173 VGND.n3172 0.40893
R6011 VGND.n1704 VGND.n1703 0.403977
R6012 VGND.n1737 VGND.n1736 0.403309
R6013 VGND.n71 VGND.n41 0.399982
R6014 VGND.n3249 VGND.n36 0.399038
R6015 VGND.n3244 VGND.n3243 0.397375
R6016 VGND.n3191 VGND.n3164 0.397302
R6017 VGND.n3191 VGND.n3158 0.395849
R6018 VGND.n2593 VGND.n954 0.394487
R6019 VGND.n3207 VGND.n80 0.392972
R6020 VGND.n70 VGND.n69 0.392942
R6021 VGND.n3207 VGND.n3150 0.391664
R6022 VGND.n69 VGND.n36 0.391488
R6023 VGND.n2349 VGND.n1027 0.389854
R6024 VGND.n2346 VGND.n2345 0.389854
R6025 VGND.n2341 VGND.n1034 0.389854
R6026 VGND.n1038 VGND.n1036 0.389854
R6027 VGND.n2232 VGND.n2220 0.389854
R6028 VGND.n2239 VGND.n2219 0.389854
R6029 VGND.n2237 VGND.n2215 0.389854
R6030 VGND.n2250 VGND.n2246 0.389854
R6031 VGND.n2263 VGND.n2262 0.389854
R6032 VGND.n2151 VGND.n2131 0.389854
R6033 VGND.n2153 VGND.n2139 0.389854
R6034 VGND.n2169 VGND.n2137 0.389854
R6035 VGND.n2731 VGND.n602 0.389854
R6036 VGND.n2737 VGND.n594 0.389854
R6037 VGND.n596 VGND.n592 0.389854
R6038 VGND.n2159 VGND.n588 0.389854
R6039 VGND.n2778 VGND.n543 0.389854
R6040 VGND.n631 VGND.n545 0.389854
R6041 VGND.n637 VGND.n629 0.389854
R6042 VGND.n634 VGND.n621 0.389854
R6043 VGND.n613 VGND.n612 0.389854
R6044 VGND.n653 VGND.n610 0.389854
R6045 VGND.n659 VGND.n658 0.389854
R6046 VGND.n2961 VGND.n2960 0.389854
R6047 VGND.n102 VGND.n35 0.388
R6048 VGND.n1739 VGND.n1738 0.388
R6049 VGND.n1737 VGND.n1065 0.388
R6050 VGND.n1543 VGND.n1304 0.385034
R6051 VGND.n3246 VGND.n3244 0.384513
R6052 VGND.n3226 VGND.n80 0.382142
R6053 VGND.n1702 VGND.n1011 0.380698
R6054 VGND.n3226 VGND.n79 0.377287
R6055 VGND VGND.n2568 0.376645
R6056 VGND.n1704 VGND.n1022 0.3725
R6057 VGND.n3203 VGND.n3150 0.371646
R6058 VGND.n1542 VGND.n1305 0.368482
R6059 VGND.n2283 VGND.n2282 0.365519
R6060 VGND.n2812 VGND.n507 0.365519
R6061 VGND.n2176 VGND.n2137 0.365519
R6062 VGND.n2135 VGND.n534 0.364266
R6063 VGND.n2179 VGND.n2178 0.364266
R6064 VGND.n2868 VGND 0.361526
R6065 VGND.n1839 VGND 0.361526
R6066 VGND.n2044 VGND 0.361526
R6067 VGND.n1589 VGND.n724 0.356056
R6068 VGND.n1586 VGND.n719 0.355071
R6069 VGND.n835 VGND.n834 0.3505
R6070 VGND.n1739 VGND.n1737 0.34884
R6071 VGND.n1703 VGND.n970 0.348815
R6072 VGND.n2351 VGND.n1022 0.341184
R6073 VGND.n3255 VGND.n26 0.337254
R6074 VGND.n2593 VGND.n2592 0.332643
R6075 VGND.n1703 VGND.n1702 0.332643
R6076 VGND.n1736 VGND.n1735 0.332643
R6077 VGND.n1226 VGND.n1225 0.327796
R6078 VGND.n3019 VGND.n291 0.3255
R6079 VGND.n3015 VGND.n305 0.3255
R6080 VGND.n3112 VGND.n3111 0.324946
R6081 VGND.n1231 VGND.n0 0.324513
R6082 VGND.n2356 VGND.n2355 0.31685
R6083 VGND.n1245 VGND.n1244 0.314886
R6084 VGND.n1239 VGND.n3 0.309856
R6085 VGND.n1570 VGND.n1010 0.309762
R6086 VGND.n1740 VGND.n1739 0.302466
R6087 VGND.n809 VGND.n310 0.3005
R6088 VGND.n3002 VGND.n3001 0.3005
R6089 VGND.n1205 VGND.n1204 0.3005
R6090 VGND.n1593 VGND.n1592 0.300032
R6091 VGND.n3230 VGND.n3229 0.299413
R6092 VGND.n1892 VGND.n1746 0.292515
R6093 VGND.n1856 VGND.n489 0.292515
R6094 VGND.n2929 VGND.n2928 0.292515
R6095 VGND.n336 VGND.n333 0.291409
R6096 VGND.n2817 VGND.n344 0.291409
R6097 VGND.n2956 VGND.n2955 0.291409
R6098 VGND.n1744 VGND.n1741 0.289991
R6099 VGND.n3247 VGND.n41 0.288821
R6100 VGND.n3247 VGND.n3246 0.287909
R6101 VGND.n3003 VGND.n3002 0.2755
R6102 VGND.n2396 VGND.n998 0.275399
R6103 VGND.n2395 VGND.n999 0.275399
R6104 VGND.n2402 VGND.n994 0.275399
R6105 VGND.n2404 VGND.n2403 0.275399
R6106 VGND.n2410 VGND.n991 0.275399
R6107 VGND.n2417 VGND.n987 0.275399
R6108 VGND.n2419 VGND.n2418 0.275399
R6109 VGND.n2692 VGND.n710 0.275399
R6110 VGND.n2691 VGND.n711 0.275399
R6111 VGND.n2687 VGND.n2686 0.275399
R6112 VGND.n1215 VGND.n1214 0.274029
R6113 VGND.n1228 VGND.n1220 0.271104
R6114 VGND.n1227 VGND.n1223 0.271104
R6115 VGND.n2332 VGND 0.268181
R6116 VGND VGND.n2138 0.268181
R6117 VGND.n647 VGND 0.268181
R6118 VGND.n1235 VGND.n1229 0.268163
R6119 VGND.n729 VGND.n726 0.26675
R6120 VGND.n2672 VGND.n721 0.266551
R6121 VGND.n3017 VGND.n299 0.262566
R6122 VGND.n2666 VGND.n2665 0.259011
R6123 VGND.n2665 VGND.n2664 0.259011
R6124 VGND.n2664 VGND.n2663 0.259011
R6125 VGND.n2663 VGND.n2662 0.259011
R6126 VGND.n753 VGND.n752 0.259011
R6127 VGND.n752 VGND.n169 0.259011
R6128 VGND.n3130 VGND.n169 0.259011
R6129 VGND.n832 VGND.n315 0.258833
R6130 VGND.n2955 VGND.n2954 0.258833
R6131 VGND.n2590 VGND.n2589 0.258833
R6132 VGND.n3282 VGND.n3281 0.258833
R6133 VGND.n1541 VGND.n1540 0.258565
R6134 VGND.n2638 VGND.n2637 0.258295
R6135 VGND.n1738 VGND.n1079 0.253965
R6136 VGND.n3233 VGND.n3232 0.253
R6137 VGND.n3248 VGND.n37 0.252092
R6138 VGND.n3249 VGND.n3248 0.251296
R6139 VGND.n3252 VGND.n3251 0.2505
R6140 VGND.n3248 VGND.n3247 0.2505
R6141 VGND.n2583 VGND.n2582 0.248699
R6142 VGND.n1211 VGND.n1210 0.245237
R6143 VGND.n1537 VGND.n1536 0.245222
R6144 VGND.n1553 VGND.n1290 0.245222
R6145 VGND.n2678 VGND.n721 0.243398
R6146 VGND.n3254 VGND.n3253 0.239337
R6147 VGND.n1592 VGND.n1591 0.238962
R6148 VGND.n2978 VGND.n333 0.238517
R6149 VGND.n1671 VGND.n1670 0.233227
R6150 VGND.n1907 VGND.n1650 0.233227
R6151 VGND.n1937 VGND.n1936 0.233227
R6152 VGND.n1260 VGND.n1173 0.233
R6153 VGND.n1234 VGND.n1233 0.232837
R6154 VGND.n75 VGND.n64 0.23175
R6155 VGND.n3125 VGND.n171 0.231578
R6156 VGND.n3001 VGND.n315 0.2255
R6157 VGND.n1574 VGND.n1002 0.223856
R6158 VGND.n2446 VGND.n971 0.223856
R6159 VGND.n3177 VGND.n83 0.22119
R6160 VGND.n40 VGND.n31 0.218488
R6161 VGND.n1239 VGND.n1238 0.216779
R6162 VGND.n1240 VGND.n1237 0.216779
R6163 VGND.n3245 VGND.n32 0.210866
R6164 VGND.n40 VGND.n39 0.205163
R6165 VGND.n39 VGND.n32 0.204516
R6166 VGND.n1155 VGND.n1150 0.203625
R6167 VGND.n85 VGND.n45 0.202674
R6168 VGND.n754 VGND.n753 0.202628
R6169 VGND.n809 VGND.n308 0.2005
R6170 VGND.n2135 VGND.n2134 0.198514
R6171 VGND.n2178 VGND.n467 0.198514
R6172 VGND.n2134 VGND.n468 0.197638
R6173 VGND.n2871 VGND.n467 0.197638
R6174 VGND.n489 VGND.n487 0.197423
R6175 VGND.n2997 VGND.n2996 0.197423
R6176 VGND.n2059 VGND.n1065 0.197423
R6177 VGND.n2928 VGND.n395 0.197423
R6178 VGND.n1743 VGND.n1742 0.194439
R6179 VGND.n744 VGND.n743 0.193248
R6180 VGND.n2870 VGND.n468 0.191226
R6181 VGND.n2177 VGND.n2135 0.190358
R6182 VGND.n992 VGND 0.189493
R6183 VGND.n832 VGND.n357 0.18703
R6184 VGND.n2954 VGND.n357 0.18703
R6185 VGND.n35 VGND.n33 0.185946
R6186 VGND.n327 VGND.n324 0.185624
R6187 VGND.n330 VGND.n328 0.185624
R6188 VGND.n730 VGND.n729 0.1855
R6189 VGND.n3250 VGND.n35 0.185359
R6190 VGND.n3152 VGND 0.18431
R6191 VGND.n3278 VGND.n9 0.181549
R6192 VGND.n1745 VGND.n1744 0.180043
R6193 VGND.n967 VGND.n714 0.17751
R6194 VGND.n2577 VGND.n963 0.17751
R6195 VGND.n2576 VGND.n964 0.17751
R6196 VGND.n2454 VGND.n2453 0.17751
R6197 VGND.n2560 VGND.n2559 0.17751
R6198 VGND.n2540 VGND.n2487 0.17751
R6199 VGND.n2539 VGND.n2536 0.17751
R6200 VGND.n2535 VGND.n2488 0.17751
R6201 VGND.n2532 VGND.n2531 0.17751
R6202 VGND.n2525 VGND.n2498 0.17751
R6203 VGND.n2524 VGND.n2522 0.17751
R6204 VGND.n2521 VGND.n2520 0.17751
R6205 VGND.n2517 VGND.n2515 0.17751
R6206 VGND.n3020 VGND.n3019 0.1755
R6207 VGND.n2871 VGND.n2870 0.173484
R6208 VGND.n3127 VGND.n168 0.171061
R6209 VGND.n2954 VGND.n2953 0.170123
R6210 VGND.n1740 VGND 0.168495
R6211 VGND.n39 VGND.n35 0.167167
R6212 VGND.n1225 VGND.n1223 0.166826
R6213 VGND.n2447 VGND.n2446 0.166571
R6214 VGND.n2178 VGND.n2177 0.165201
R6215 VGND.n833 VGND.n832 0.165134
R6216 VGND VGND.n2867 0.164603
R6217 VGND.n1816 VGND 0.164603
R6218 VGND VGND.n2043 0.164603
R6219 VGND.n1539 VGND.n10 0.162882
R6220 VGND.n2447 VGND.n970 0.161835
R6221 VGND.n2587 VGND.n954 0.159519
R6222 VGND.n3277 VGND 0.159365
R6223 VGND.n1538 VGND.n1306 0.159008
R6224 VGND.n3196 VGND.n3195 0.158313
R6225 VGND.n3161 VGND.n3151 0.158313
R6226 VGND.n3179 VGND.n3174 0.158313
R6227 VGND.n2645 VGND.n733 0.158127
R6228 VGND.n940 VGND.n734 0.158127
R6229 VGND.n735 VGND.n175 0.158127
R6230 VGND.n737 VGND.n736 0.158127
R6231 VGND.n748 VGND.n747 0.158127
R6232 VGND.n773 VGND.n732 0.158127
R6233 VGND.n2625 VGND.n731 0.158127
R6234 VGND.n751 VGND.n191 0.158127
R6235 VGND.n3132 VGND.n3131 0.158127
R6236 VGND.n1595 VGND.n1594 0.1555
R6237 VGND.n3161 VGND.n3160 0.153625
R6238 VGND.n3180 VGND.n3179 0.153625
R6239 VGND.n1156 VGND.n1092 0.153488
R6240 VGND.n1252 VGND.n1177 0.152595
R6241 VGND.n1209 VGND.n1208 0.151324
R6242 VGND.n3256 VGND.n29 0.1505
R6243 VGND.n1414 VGND.n1413 0.147888
R6244 VGND.n2960 VGND.n351 0.146508
R6245 VGND.n724 VGND.n723 0.145813
R6246 VGND.n1585 VGND.n1579 0.145813
R6247 VGND.n2570 VGND.n968 0.14432
R6248 VGND.n8 VGND 0.143615
R6249 VGND.n2640 VGND.n2639 0.142439
R6250 VGND.n738 VGND.n173 0.142439
R6251 VGND.n750 VGND.n749 0.142439
R6252 VGND.n749 VGND.n168 0.142439
R6253 VGND.n2639 VGND.n2638 0.140273
R6254 VGND.n1238 VGND.n5 0.140064
R6255 VGND.n2671 VGND.n2670 0.139306
R6256 VGND.n744 VGND.n738 0.138643
R6257 VGND.n3197 VGND.n3194 0.138
R6258 VGND.n1254 VGND.n1253 0.133357
R6259 VGND.n3256 VGND.n3255 0.132853
R6260 VGND.n874 VGND.n355 0.132731
R6261 VGND.n2567 VGND.n2448 0.131237
R6262 VGND.n1234 VGND.n0 0.13045
R6263 VGND.n833 VGND.n831 0.129935
R6264 VGND.n834 VGND.n833 0.129667
R6265 VGND.n1223 VGND.n1220 0.127728
R6266 VGND.n2643 VGND.n2642 0.126668
R6267 VGND.n1540 VGND.n1272 0.126176
R6268 VGND.n121 VGND.n30 0.126163
R6269 VGND.n3075 VGND.n224 0.123973
R6270 VGND.n73 VGND.n58 0.122868
R6271 VGND.n2641 VGND.n172 0.122579
R6272 VGND.n3279 VGND.n3278 0.122286
R6273 VGND.n2570 VGND 0.122194
R6274 VGND VGND.n2489 0.122194
R6275 VGND.n2226 VGND 0.122173
R6276 VGND.n2144 VGND 0.122173
R6277 VGND VGND.n646 0.122173
R6278 VGND.n3242 VGND.n3241 0.121279
R6279 VGND.n1235 VGND.n1234 0.120302
R6280 VGND.n2953 VGND.n2952 0.119731
R6281 VGND.n2675 VGND.n724 0.119019
R6282 VGND.n3225 VGND.n81 0.119019
R6283 VGND.n2449 VGND.n358 0.115799
R6284 VGND.n3124 VGND.n172 0.113818
R6285 VGND.n357 VGND.n333 0.111214
R6286 VGND.n3281 VGND.n3280 0.108503
R6287 VGND.n1544 VGND.n1303 0.106901
R6288 VGND.n3229 VGND.n3228 0.105176
R6289 VGND.n2283 VGND.n467 0.103833
R6290 VGND.n2134 VGND.n507 0.103833
R6291 VGND.n3231 VGND.n76 0.103014
R6292 VGND.n3163 VGND.n3162 0.101587
R6293 VGND.n3178 VGND.n3177 0.101587
R6294 VGND.n2284 VGND.n2283 0.0978384
R6295 VGND.n507 VGND.n506 0.0978384
R6296 VGND.n1241 VGND.n1240 0.09425
R6297 VGND.n3171 VGND.n3168 0.0939307
R6298 VGND.n894 VGND.n274 0.0935
R6299 VGND.n1216 VGND.n1215 0.0883906
R6300 VGND.n45 VGND.n44 0.0870385
R6301 VGND.n2411 VGND 0.086406
R6302 VGND.n1744 VGND.n1743 0.0806724
R6303 VGND.n1256 VGND.n1175 0.0806724
R6304 VGND.n2971 VGND.n339 0.0798388
R6305 VGND.t109 VGND.t93 0.0785455
R6306 VGND.n1415 VGND.n1378 0.0783116
R6307 VGND.n1898 VGND.n1650 0.0780758
R6308 VGND.n1936 VGND.n1627 0.0780758
R6309 VGND.n2177 VGND.n2176 0.078
R6310 VGND.n2514 VGND.n2500 0.0770894
R6311 VGND.n2870 VGND.n2869 0.0755
R6312 VGND.n2996 VGND.n315 0.0755
R6313 VGND.n3285 VGND.n3284 0.0755
R6314 VGND.n3254 VGND.n30 0.0736479
R6315 VGND.n3040 VGND 0.0714541
R6316 VGND.n3217 VGND.n63 0.0701203
R6317 VGND.n1182 VGND.n1177 0.0688498
R6318 VGND.n1243 VGND.n1220 0.0685693
R6319 VGND.n1153 VGND.n1152 0.0664574
R6320 VGND.n3044 VGND.n3043 0.0664574
R6321 VGND.n2953 VGND.n358 0.0661874
R6322 VGND.n2928 VGND.n394 0.066141
R6323 VGND.n1852 VGND.n489 0.066141
R6324 VGND.n1209 VGND.n1187 0.0658846
R6325 VGND.n1241 VGND.n1235 0.065599
R6326 VGND.n1257 VGND.n1256 0.0646604
R6327 VGND.n2358 VGND.n2357 0.0638663
R6328 VGND.n2365 VGND.n1014 0.0638663
R6329 VGND.n2364 VGND.n1012 0.0638663
R6330 VGND.n2371 VGND.n1011 0.0638663
R6331 VGND.n2374 VGND.n2373 0.0638663
R6332 VGND.n2381 VGND.n1007 0.0638663
R6333 VGND.n2380 VGND.n1005 0.0638663
R6334 VGND.n1004 VGND.n1001 0.0638663
R6335 VGND.n2389 VGND.n2388 0.0638663
R6336 VGND.n1969 VGND.n1081 0.0638663
R6337 VGND.n1975 VGND.n1973 0.0638663
R6338 VGND.n1974 VGND.n1077 0.0638663
R6339 VGND.n1982 VGND.n1981 0.0638663
R6340 VGND.n1075 VGND.n1074 0.0638663
R6341 VGND.n1990 VGND.n1988 0.0638663
R6342 VGND.n1989 VGND.n1072 0.0638663
R6343 VGND.n2000 VGND.n1999 0.0638663
R6344 VGND.n1070 VGND.n1064 0.0638663
R6345 VGND.n1059 VGND.n1056 0.0638663
R6346 VGND.n2325 VGND.n2324 0.0638663
R6347 VGND.n1705 VGND.n1057 0.0638663
R6348 VGND.n1734 VGND.n1706 0.0638663
R6349 VGND.n1731 VGND.n1730 0.0638663
R6350 VGND.n1726 VGND.n1708 0.0638663
R6351 VGND.n1725 VGND.n1722 0.0638663
R6352 VGND.n1721 VGND.n1717 0.0638663
R6353 VGND.n1718 VGND.n1016 0.0638663
R6354 VGND.n1191 VGND.n1179 0.063
R6355 VGND.n1149 VGND.n266 0.0611996
R6356 VGND.n1218 VGND.n1217 0.0603131
R6357 VGND.n1238 VGND.n1237 0.0603131
R6358 VGND.n1183 VGND.n1182 0.0601154
R6359 VGND.n1206 VGND.n1205 0.0597352
R6360 VGND.n1208 VGND.n1189 0.0593608
R6361 VGND.n1249 VGND.n1248 0.0558571
R6362 VGND VGND.n2569 0.0558155
R6363 VGND.n2495 VGND 0.0558155
R6364 VGND.n170 VGND.n156 0.0530424
R6365 VGND.n73 VGND.n72 0.0528256
R6366 VGND.n3243 VGND.n3242 0.0528256
R6367 VGND.n2446 VGND.n2445 0.0520436
R6368 VGND.n3253 VGND.n3252 0.0515
R6369 VGND.n1415 VGND.n1414 0.0510435
R6370 VGND.n1233 VGND.n1232 0.0509808
R6371 VGND.n834 VGND.n828 0.0505
R6372 VGND.n1261 VGND.n1 0.0505
R6373 VGND.n1584 VGND.n1583 0.0489375
R6374 VGND.n2662 VGND.n2661 0.0489043
R6375 VGND.n2448 VGND.n2447 0.0474402
R6376 VGND.n1408 VGND.n1273 0.0460882
R6377 VGND.n3179 VGND.n3178 0.0446176
R6378 VGND.n3163 VGND.n3161 0.0446176
R6379 VGND.n3196 VGND.n3153 0.0446176
R6380 VGND.n1583 VGND.n1579 0.0443356
R6381 VGND.n2661 VGND.n2660 0.044162
R6382 VGND.n1236 VGND.n1219 0.0437558
R6383 VGND.n3129 VGND.n170 0.0434537
R6384 VGND.n112 VGND.n97 0.0430249
R6385 VGND VGND.n3288 0.0416676
R6386 VGND.n2644 VGND.n2643 0.0416504
R6387 VGND.n1236 VGND.n1218 0.0403754
R6388 VGND.n3274 VGND.n3273 0.0399068
R6389 VGND.n270 VGND.t87 0.0364339
R6390 VGND.n3276 VGND.n3275 0.0345909
R6391 VGND.n1535 VGND.n1306 0.0338333
R6392 VGND.n2867 VGND 0.0333205
R6393 VGND.n1816 VGND 0.0333205
R6394 VGND.n2043 VGND 0.0333205
R6395 VGND.n3036 VGND.n3035 0.0332465
R6396 VGND.n831 VGND.n275 0.0332051
R6397 VGND.n3288 VGND.n0 0.0316881
R6398 VGND.n2636 VGND.n777 0.029221
R6399 VGND.n3124 VGND.n173 0.0291215
R6400 VGND.n1412 VGND.n1411 0.0288912
R6401 VGND.n268 VGND.n266 0.0288019
R6402 VGND.n1151 VGND.n273 0.0288019
R6403 VGND.n2637 VGND.n2636 0.0286818
R6404 VGND.n777 VGND.n776 0.0286818
R6405 VGND.n3286 VGND.n2 0.0282356
R6406 VGND.n1262 VGND.n1261 0.0280862
R6407 VGND.n1260 VGND.n1259 0.0280862
R6408 VGND.n1262 VGND.n1174 0.0272241
R6409 VGND.n2635 VGND.n778 0.0266759
R6410 VGND.n1249 VGND.n1180 0.0260682
R6411 VGND.n1251 VGND.n1178 0.0252302
R6412 VGND.n1893 VGND.n1892 0.0248346
R6413 VGND.n1888 VGND.n1758 0.0248346
R6414 VGND.n1762 VGND.n1761 0.0248346
R6415 VGND.n1883 VGND.n1763 0.0248346
R6416 VGND.n1879 VGND.n1878 0.0248346
R6417 VGND.n1874 VGND.n1778 0.0248346
R6418 VGND.n1782 VGND.n1781 0.0248346
R6419 VGND.n1869 VGND.n1783 0.0248346
R6420 VGND.n1865 VGND.n1864 0.0248346
R6421 VGND.n2256 VGND.n692 0.0248346
R6422 VGND.n2707 VGND.n694 0.0248346
R6423 VGND.n2200 VGND.n2199 0.0248346
R6424 VGND.n2197 VGND.n2185 0.0248346
R6425 VGND.n2206 VGND.n2196 0.0248346
R6426 VGND.n2193 VGND.n2190 0.0248346
R6427 VGND.n2429 VGND.n2428 0.0248346
R6428 VGND.n980 VGND.n979 0.0248346
R6429 VGND.n2436 VGND.n2435 0.0248346
R6430 VGND.n2292 VGND.n2072 0.0248346
R6431 VGND.n2288 VGND.n2077 0.0248346
R6432 VGND.n2080 VGND.n2079 0.0248346
R6433 VGND.n2282 VGND.n2081 0.0248346
R6434 VGND.n2278 VGND.n2277 0.0248346
R6435 VGND.n2273 VGND.n2120 0.0248346
R6436 VGND.n2126 VGND.n2123 0.0248346
R6437 VGND.n2268 VGND.n2127 0.0248346
R6438 VGND.n2717 VGND.n685 0.0248346
R6439 VGND.n2846 VGND.n497 0.0248346
R6440 VGND.n503 VGND.n500 0.0248346
R6441 VGND.n2840 VGND.n504 0.0248346
R6442 VGND.n2812 VGND.n2811 0.0248346
R6443 VGND.n2805 VGND.n514 0.0248346
R6444 VGND.n521 VGND.n517 0.0248346
R6445 VGND.n2799 VGND.n522 0.0248346
R6446 VGND.n2793 VGND.n2792 0.0248346
R6447 VGND.n2786 VGND.n531 0.0248346
R6448 VGND.n2772 VGND.n2771 0.0248346
R6449 VGND.n2768 VGND.n571 0.0248346
R6450 VGND.n2752 VGND.n574 0.0248346
R6451 VGND.n2758 VGND.n578 0.0248346
R6452 VGND.n2761 VGND.n2757 0.0248346
R6453 VGND.n2472 VGND.n2470 0.0248346
R6454 VGND.n2477 VGND.n2462 0.0248346
R6455 VGND.n2466 VGND.n2450 0.0248346
R6456 VGND.n2550 VGND.n2451 0.0248346
R6457 VGND VGND.n2226 0.0248346
R6458 VGND.n2144 VGND 0.0248346
R6459 VGND.n646 VGND 0.0248346
R6460 VGND.n2913 VGND.n2912 0.0248346
R6461 VGND.n2908 VGND.n437 0.0248346
R6462 VGND.n450 VGND.n440 0.0248346
R6463 VGND.n447 VGND.n446 0.0248346
R6464 VGND.n2901 VGND.n448 0.0248346
R6465 VGND.n2898 VGND.n2897 0.0248346
R6466 VGND.n2890 VGND.n459 0.0248346
R6467 VGND.n2878 VGND.n463 0.0248346
R6468 VGND.n2884 VGND.n2882 0.0248346
R6469 VGND.n1251 VGND.n1250 0.0244362
R6470 VGND.n11 VGND.n10 0.0221346
R6471 VGND.n1237 VGND.n1236 0.0204377
R6472 VGND.n2642 VGND.n2641 0.0203598
R6473 VGND.n1154 VGND.n1153 0.0193442
R6474 VGND.n1242 VGND.n1219 0.01925
R6475 VGND.n1156 VGND.n1155 0.0189524
R6476 VGND.t108 VGND.n270 0.0180899
R6477 VGND.n2411 VGND 0.0176812
R6478 VGND.n3199 VGND.n3198 0.0173018
R6479 VGND.n2643 VGND.n2640 0.016271
R6480 VGND.n3197 VGND.n3196 0.016125
R6481 VGND.n1410 VGND.n1409 0.0153026
R6482 VGND.n267 VGND.n224 0.0143393
R6483 VGND.n3233 VGND.n75 0.01425
R6484 VGND.n3287 VGND.n3286 0.0135435
R6485 VGND.n1410 VGND.n1408 0.0119353
R6486 VGND.n270 VGND.n269 0.0115828
R6487 VGND.n2569 VGND 0.0115631
R6488 VGND VGND.n2495 0.0115631
R6489 VGND.n74 VGND.n60 0.00861884
R6490 VGND.n2661 VGND.n754 0.00847872
R6491 VGND.n2588 VGND.n2587 0.00838733
R6492 VGND.n3234 VGND.n60 0.00831506
R6493 VGND.n1207 VGND.n7 0.00764286
R6494 VGND.n1584 VGND.n1581 0.00739338
R6495 VGND.n2641 VGND.n171 0.00725676
R6496 VGND.n3042 VGND.n3041 0.00645238
R6497 VGND.n3216 VGND.n79 0.0055975
R6498 VGND.n750 VGND.n744 0.00429673
R6499 VGND.n1539 VGND.n1538 0.00297529
R6500 VGND.n3275 VGND.n3274 0.00236567
R6501 VGND.n269 VGND.t0 0.00163108
R6502 VGND.n2676 VGND.n723 0.00154167
R6503 VGND.n2637 VGND.n776 0.00142822
R6504 VGND.n3042 VGND.n267 0.00140909
R6505 VGND.n3231 VGND.n3230 0.00139297
R6506 VGND.n269 VGND.t102 0.00136679
R6507 VGND.n1261 VGND.n1260 0.00136207
R6508 VGND.n1240 VGND.n1239 0.00125453
R6509 VGND.n1153 VGND.n1151 0.00112814
R6510 VGND.n3199 VGND.n3153 0.0011252
R6511 VGND.n3043 VGND.n266 0.0010144
R6512 VGND.n1244 VGND.n1219 0.00100302
R6513 VGND.n1243 VGND.n1242 0.00099505
R6514 VGND.n1250 VGND.n1249 0.000973485
R6515 VGND.n1585 VGND.n1584 0.000959559
R6516 VGND.n1240 VGND.n1219 0.000751509
R6517 VGND.n1242 VGND.n1241 0.000747525
R6518 VGND.n1306 VGND.n11 0.000612309
R6519 ua[5].t1 ua[5].t0 359.057
R6520 ua[5] ua[5].t1 244.087
R6521 a_16597_7688.n93 a_16597_7688.t8 669.811
R6522 a_16597_7688.t8 a_16597_7688.n92 669.811
R6523 a_16597_7688.t10 a_16597_7688.n18 669.811
R6524 a_16597_7688.n91 a_16597_7688.t10 669.811
R6525 a_16597_7688.t36 a_16597_7688.n88 669.811
R6526 a_16597_7688.n89 a_16597_7688.t36 669.811
R6527 a_16597_7688.n86 a_16597_7688.t4 669.811
R6528 a_16597_7688.t4 a_16597_7688.n21 669.811
R6529 a_16597_7688.n84 a_16597_7688.t24 669.811
R6530 a_16597_7688.t24 a_16597_7688.n83 669.811
R6531 a_16597_7688.t38 a_16597_7688.n22 669.811
R6532 a_16597_7688.n79 a_16597_7688.t38 669.811
R6533 a_16597_7688.t18 a_16597_7688.n76 669.811
R6534 a_16597_7688.n77 a_16597_7688.t18 669.811
R6535 a_16597_7688.n74 a_16597_7688.t28 669.811
R6536 a_16597_7688.t28 a_16597_7688.n25 669.811
R6537 a_16597_7688.n72 a_16597_7688.t32 669.811
R6538 a_16597_7688.t32 a_16597_7688.n71 669.811
R6539 a_16597_7688.t30 a_16597_7688.n26 669.811
R6540 a_16597_7688.n67 a_16597_7688.t30 669.811
R6541 a_16597_7688.t26 a_16597_7688.n64 669.811
R6542 a_16597_7688.n65 a_16597_7688.t26 669.811
R6543 a_16597_7688.n62 a_16597_7688.t2 669.811
R6544 a_16597_7688.t2 a_16597_7688.n29 669.811
R6545 a_16597_7688.n60 a_16597_7688.t22 669.811
R6546 a_16597_7688.t22 a_16597_7688.n59 669.811
R6547 a_16597_7688.t16 a_16597_7688.n30 669.811
R6548 a_16597_7688.n55 a_16597_7688.t16 669.811
R6549 a_16597_7688.t14 a_16597_7688.n52 669.811
R6550 a_16597_7688.n53 a_16597_7688.t14 669.811
R6551 a_16597_7688.n50 a_16597_7688.t12 669.811
R6552 a_16597_7688.t12 a_16597_7688.n33 669.811
R6553 a_16597_7688.n48 a_16597_7688.t20 669.811
R6554 a_16597_7688.t20 a_16597_7688.n47 669.811
R6555 a_16597_7688.t34 a_16597_7688.n34 669.811
R6556 a_16597_7688.n43 a_16597_7688.t34 669.811
R6557 a_16597_7688.t6 a_16597_7688.n40 669.811
R6558 a_16597_7688.n41 a_16597_7688.t6 669.811
R6559 a_16597_7688.n38 a_16597_7688.t0 669.811
R6560 a_16597_7688.t0 a_16597_7688.n37 669.811
R6561 a_16597_7688.t42 a_16597_7688.n3 669.811
R6562 a_16597_7688.n4 a_16597_7688.t42 669.811
R6563 a_16597_7688.n6 a_16597_7688.t40 669.811
R6564 a_16597_7688.t40 a_16597_7688.n5 669.811
R6565 a_16597_7688.n95 a_16597_7688.t44 86.5538
R6566 a_16597_7688.n17 a_16597_7688.t9 8.37725
R6567 a_16597_7688.n2 a_16597_7688.t41 8.37725
R6568 a_16597_7688.n36 a_16597_7688.n35 6.72425
R6569 a_16597_7688.n45 a_16597_7688.n44 6.72425
R6570 a_16597_7688.n32 a_16597_7688.n31 6.72425
R6571 a_16597_7688.n57 a_16597_7688.n56 6.72425
R6572 a_16597_7688.n28 a_16597_7688.n27 6.72425
R6573 a_16597_7688.n69 a_16597_7688.n68 6.72425
R6574 a_16597_7688.n24 a_16597_7688.n23 6.72425
R6575 a_16597_7688.n81 a_16597_7688.n80 6.72425
R6576 a_16597_7688.n20 a_16597_7688.n19 6.72425
R6577 a_16597_7688.n108 a_16597_7688.n107 6.72425
R6578 a_16597_7688.n5 a_16597_7688.n2 3.01952
R6579 a_16597_7688.n92 a_16597_7688.n17 3.01952
R6580 a_16597_7688.n42 a_16597_7688.n36 2.80485
R6581 a_16597_7688.n46 a_16597_7688.n45 2.80485
R6582 a_16597_7688.n54 a_16597_7688.n32 2.80485
R6583 a_16597_7688.n58 a_16597_7688.n57 2.80485
R6584 a_16597_7688.n66 a_16597_7688.n28 2.80485
R6585 a_16597_7688.n70 a_16597_7688.n69 2.80485
R6586 a_16597_7688.n78 a_16597_7688.n24 2.80485
R6587 a_16597_7688.n82 a_16597_7688.n81 2.80485
R6588 a_16597_7688.n90 a_16597_7688.n20 2.80485
R6589 a_16597_7688.n107 a_16597_7688.n0 2.80485
R6590 a_16597_7688.n36 a_16597_7688.n8 1.94555
R6591 a_16597_7688.n45 a_16597_7688.n9 1.94555
R6592 a_16597_7688.n32 a_16597_7688.n10 1.94555
R6593 a_16597_7688.n57 a_16597_7688.n11 1.94555
R6594 a_16597_7688.n28 a_16597_7688.n12 1.94555
R6595 a_16597_7688.n69 a_16597_7688.n13 1.94555
R6596 a_16597_7688.n24 a_16597_7688.n14 1.94555
R6597 a_16597_7688.n81 a_16597_7688.n15 1.94555
R6598 a_16597_7688.n20 a_16597_7688.n16 1.94555
R6599 a_16597_7688.n7 a_16597_7688.n2 1.94555
R6600 a_16597_7688.n94 a_16597_7688.n17 1.94555
R6601 a_16597_7688.n107 a_16597_7688.n106 1.94555
R6602 a_16597_7688.n35 a_16597_7688.t7 1.6535
R6603 a_16597_7688.n35 a_16597_7688.t35 1.6535
R6604 a_16597_7688.n44 a_16597_7688.t21 1.6535
R6605 a_16597_7688.n44 a_16597_7688.t13 1.6535
R6606 a_16597_7688.n31 a_16597_7688.t15 1.6535
R6607 a_16597_7688.n31 a_16597_7688.t17 1.6535
R6608 a_16597_7688.n56 a_16597_7688.t23 1.6535
R6609 a_16597_7688.n56 a_16597_7688.t3 1.6535
R6610 a_16597_7688.n27 a_16597_7688.t27 1.6535
R6611 a_16597_7688.n27 a_16597_7688.t31 1.6535
R6612 a_16597_7688.n68 a_16597_7688.t33 1.6535
R6613 a_16597_7688.n68 a_16597_7688.t29 1.6535
R6614 a_16597_7688.n23 a_16597_7688.t19 1.6535
R6615 a_16597_7688.n23 a_16597_7688.t39 1.6535
R6616 a_16597_7688.n80 a_16597_7688.t25 1.6535
R6617 a_16597_7688.n80 a_16597_7688.t5 1.6535
R6618 a_16597_7688.n19 a_16597_7688.t37 1.6535
R6619 a_16597_7688.n19 a_16597_7688.t11 1.6535
R6620 a_16597_7688.n108 a_16597_7688.t43 1.6535
R6621 a_16597_7688.t1 a_16597_7688.n108 1.6535
R6622 a_16597_7688.n105 a_16597_7688.n7 1.21883
R6623 a_16597_7688.n106 a_16597_7688.n105 0.928385
R6624 a_16597_7688.n104 a_16597_7688.n8 0.928385
R6625 a_16597_7688.n103 a_16597_7688.n9 0.928385
R6626 a_16597_7688.n102 a_16597_7688.n10 0.928385
R6627 a_16597_7688.n101 a_16597_7688.n11 0.928385
R6628 a_16597_7688.n100 a_16597_7688.n12 0.928385
R6629 a_16597_7688.n99 a_16597_7688.n13 0.928385
R6630 a_16597_7688.n98 a_16597_7688.n14 0.928385
R6631 a_16597_7688.n97 a_16597_7688.n15 0.928385
R6632 a_16597_7688.n96 a_16597_7688.n16 0.928385
R6633 a_16597_7688.n95 a_16597_7688.n94 0.928385
R6634 a_16597_7688.n7 a_16597_7688.n6 0.681961
R6635 a_16597_7688.n94 a_16597_7688.n93 0.681961
R6636 a_16597_7688.n39 a_16597_7688.n8 0.467287
R6637 a_16597_7688.n49 a_16597_7688.n9 0.467287
R6638 a_16597_7688.n51 a_16597_7688.n10 0.467287
R6639 a_16597_7688.n61 a_16597_7688.n11 0.467287
R6640 a_16597_7688.n63 a_16597_7688.n12 0.467287
R6641 a_16597_7688.n73 a_16597_7688.n13 0.467287
R6642 a_16597_7688.n75 a_16597_7688.n14 0.467287
R6643 a_16597_7688.n85 a_16597_7688.n15 0.467287
R6644 a_16597_7688.n87 a_16597_7688.n16 0.467287
R6645 a_16597_7688.n106 a_16597_7688.n1 0.467287
R6646 a_16597_7688.n5 a_16597_7688.n4 0.429848
R6647 a_16597_7688.n41 a_16597_7688.n37 0.429848
R6648 a_16597_7688.n47 a_16597_7688.n43 0.429848
R6649 a_16597_7688.n53 a_16597_7688.n33 0.429848
R6650 a_16597_7688.n59 a_16597_7688.n55 0.429848
R6651 a_16597_7688.n65 a_16597_7688.n29 0.429848
R6652 a_16597_7688.n71 a_16597_7688.n67 0.429848
R6653 a_16597_7688.n77 a_16597_7688.n25 0.429848
R6654 a_16597_7688.n83 a_16597_7688.n79 0.429848
R6655 a_16597_7688.n89 a_16597_7688.n21 0.429848
R6656 a_16597_7688.n92 a_16597_7688.n91 0.429848
R6657 a_16597_7688.n6 a_16597_7688.n3 0.429848
R6658 a_16597_7688.n40 a_16597_7688.n38 0.429848
R6659 a_16597_7688.n48 a_16597_7688.n34 0.429848
R6660 a_16597_7688.n52 a_16597_7688.n50 0.429848
R6661 a_16597_7688.n60 a_16597_7688.n30 0.429848
R6662 a_16597_7688.n64 a_16597_7688.n62 0.429848
R6663 a_16597_7688.n72 a_16597_7688.n26 0.429848
R6664 a_16597_7688.n76 a_16597_7688.n74 0.429848
R6665 a_16597_7688.n84 a_16597_7688.n22 0.429848
R6666 a_16597_7688.n88 a_16597_7688.n86 0.429848
R6667 a_16597_7688.n93 a_16597_7688.n18 0.429848
R6668 a_16597_7688.n105 a_16597_7688.n104 0.290941
R6669 a_16597_7688.n104 a_16597_7688.n103 0.290941
R6670 a_16597_7688.n103 a_16597_7688.n102 0.290941
R6671 a_16597_7688.n102 a_16597_7688.n101 0.290941
R6672 a_16597_7688.n101 a_16597_7688.n100 0.290941
R6673 a_16597_7688.n100 a_16597_7688.n99 0.290941
R6674 a_16597_7688.n99 a_16597_7688.n98 0.290941
R6675 a_16597_7688.n98 a_16597_7688.n97 0.290941
R6676 a_16597_7688.n97 a_16597_7688.n96 0.290941
R6677 a_16597_7688.n96 a_16597_7688.n95 0.290941
R6678 a_16597_7688.n4 a_16597_7688.n0 0.215174
R6679 a_16597_7688.n37 a_16597_7688.n0 0.215174
R6680 a_16597_7688.n42 a_16597_7688.n41 0.215174
R6681 a_16597_7688.n43 a_16597_7688.n42 0.215174
R6682 a_16597_7688.n47 a_16597_7688.n46 0.215174
R6683 a_16597_7688.n46 a_16597_7688.n33 0.215174
R6684 a_16597_7688.n54 a_16597_7688.n53 0.215174
R6685 a_16597_7688.n55 a_16597_7688.n54 0.215174
R6686 a_16597_7688.n59 a_16597_7688.n58 0.215174
R6687 a_16597_7688.n58 a_16597_7688.n29 0.215174
R6688 a_16597_7688.n66 a_16597_7688.n65 0.215174
R6689 a_16597_7688.n67 a_16597_7688.n66 0.215174
R6690 a_16597_7688.n71 a_16597_7688.n70 0.215174
R6691 a_16597_7688.n70 a_16597_7688.n25 0.215174
R6692 a_16597_7688.n78 a_16597_7688.n77 0.215174
R6693 a_16597_7688.n79 a_16597_7688.n78 0.215174
R6694 a_16597_7688.n83 a_16597_7688.n82 0.215174
R6695 a_16597_7688.n82 a_16597_7688.n21 0.215174
R6696 a_16597_7688.n90 a_16597_7688.n89 0.215174
R6697 a_16597_7688.n91 a_16597_7688.n90 0.215174
R6698 a_16597_7688.n3 a_16597_7688.n1 0.215174
R6699 a_16597_7688.n38 a_16597_7688.n1 0.215174
R6700 a_16597_7688.n40 a_16597_7688.n39 0.215174
R6701 a_16597_7688.n39 a_16597_7688.n34 0.215174
R6702 a_16597_7688.n49 a_16597_7688.n48 0.215174
R6703 a_16597_7688.n50 a_16597_7688.n49 0.215174
R6704 a_16597_7688.n52 a_16597_7688.n51 0.215174
R6705 a_16597_7688.n51 a_16597_7688.n30 0.215174
R6706 a_16597_7688.n61 a_16597_7688.n60 0.215174
R6707 a_16597_7688.n62 a_16597_7688.n61 0.215174
R6708 a_16597_7688.n64 a_16597_7688.n63 0.215174
R6709 a_16597_7688.n63 a_16597_7688.n26 0.215174
R6710 a_16597_7688.n73 a_16597_7688.n72 0.215174
R6711 a_16597_7688.n74 a_16597_7688.n73 0.215174
R6712 a_16597_7688.n76 a_16597_7688.n75 0.215174
R6713 a_16597_7688.n75 a_16597_7688.n22 0.215174
R6714 a_16597_7688.n85 a_16597_7688.n84 0.215174
R6715 a_16597_7688.n86 a_16597_7688.n85 0.215174
R6716 a_16597_7688.n88 a_16597_7688.n87 0.215174
R6717 a_16597_7688.n87 a_16597_7688.n18 0.215174
R6718 Timming_0.Vd.n1 Timming_0.Vd.t26 238.796
R6719 Timming_0.Vd.n3 Timming_0.Vd.t24 232.821
R6720 Timming_0.Vd.n1 Timming_0.Vd.t27 121.04
R6721 Timming_0.Vd.n0 Timming_0.Vd.t1 89.1547
R6722 Timming_0.Vd.n0 Timming_0.Vd.t25 87.4384
R6723 Timming_0.Vd.n19 Timming_0.Vd.n10 9.5975
R6724 Timming_0.Vd.n15 Timming_0.Vd.n14 9.59719
R6725 Timming_0.Vd.n16 Timming_0.Vd.n13 9.59719
R6726 Timming_0.Vd.n17 Timming_0.Vd.n12 9.59719
R6727 Timming_0.Vd.n18 Timming_0.Vd.n11 9.59719
R6728 Timming_0.Vd.n20 Timming_0.Vd.n9 9.59719
R6729 Timming_0.Vd.n21 Timming_0.Vd.n8 9.59719
R6730 Timming_0.Vd.n22 Timming_0.Vd.n7 9.59719
R6731 Timming_0.Vd.n23 Timming_0.Vd.n6 9.59719
R6732 Timming_0.Vd.n24 Timming_0.Vd.n5 9.59719
R6733 Timming_0.Vd.n25 Timming_0.Vd.n4 9.59719
R6734 Timming_0.Vd.n15 Timming_0.Vd.t0 6.6127
R6735 Timming_0.Vd.n2 Timming_0.Vd.n1 5.50134
R6736 Timming_0.Vd.n10 Timming_0.Vd.t9 1.6535
R6737 Timming_0.Vd.n10 Timming_0.Vd.t6 1.6535
R6738 Timming_0.Vd.n14 Timming_0.Vd.t7 1.6535
R6739 Timming_0.Vd.n14 Timming_0.Vd.t13 1.6535
R6740 Timming_0.Vd.n13 Timming_0.Vd.t14 1.6535
R6741 Timming_0.Vd.n13 Timming_0.Vd.t20 1.6535
R6742 Timming_0.Vd.n12 Timming_0.Vd.t21 1.6535
R6743 Timming_0.Vd.n12 Timming_0.Vd.t2 1.6535
R6744 Timming_0.Vd.n11 Timming_0.Vd.t4 1.6535
R6745 Timming_0.Vd.n11 Timming_0.Vd.t16 1.6535
R6746 Timming_0.Vd.n9 Timming_0.Vd.t18 1.6535
R6747 Timming_0.Vd.n9 Timming_0.Vd.t5 1.6535
R6748 Timming_0.Vd.n8 Timming_0.Vd.t12 1.6535
R6749 Timming_0.Vd.n8 Timming_0.Vd.t10 1.6535
R6750 Timming_0.Vd.n7 Timming_0.Vd.t11 1.6535
R6751 Timming_0.Vd.n7 Timming_0.Vd.t23 1.6535
R6752 Timming_0.Vd.n6 Timming_0.Vd.t19 1.6535
R6753 Timming_0.Vd.n6 Timming_0.Vd.t22 1.6535
R6754 Timming_0.Vd.n5 Timming_0.Vd.t8 1.6535
R6755 Timming_0.Vd.n5 Timming_0.Vd.t15 1.6535
R6756 Timming_0.Vd.n4 Timming_0.Vd.t17 1.6535
R6757 Timming_0.Vd.n4 Timming_0.Vd.t3 1.6535
R6758 Timming_0.Vd.n2 Timming_0.Vd.n0 1.55579
R6759 Timming_0.Vd Timming_0.Vd.n3 0.565315
R6760 Timming_0.Vd Timming_0.Vd.n25 0.559324
R6761 Timming_0.Vd.n3 Timming_0.Vd.n2 0.315315
R6762 Timming_0.Vd.n25 Timming_0.Vd.n24 0.290941
R6763 Timming_0.Vd.n24 Timming_0.Vd.n23 0.290941
R6764 Timming_0.Vd.n23 Timming_0.Vd.n22 0.290941
R6765 Timming_0.Vd.n22 Timming_0.Vd.n21 0.290941
R6766 Timming_0.Vd.n21 Timming_0.Vd.n20 0.290941
R6767 Timming_0.Vd.n20 Timming_0.Vd.n19 0.290941
R6768 Timming_0.Vd.n19 Timming_0.Vd.n18 0.290941
R6769 Timming_0.Vd.n18 Timming_0.Vd.n17 0.290941
R6770 Timming_0.Vd.n17 Timming_0.Vd.n16 0.290941
R6771 Timming_0.Vd.n16 Timming_0.Vd.n15 0.290941
R6772 ua[2].n7 ua[2].t6 214.405
R6773 ua[2].t6 ua[2].n6 214.405
R6774 ua[2].n5 ua[2].t5 107.21
R6775 ua[2].n25 ua[2].t10 106.907
R6776 ua[2].n21 ua[2].t11 106.907
R6777 ua[2].n16 ua[2].t2 106.907
R6778 ua[2].n11 ua[2].t8 106.907
R6779 ua[2].n8 ua[2].t7 106.907
R6780 ua[2].n13 ua[2].t4 106.907
R6781 ua[2].n18 ua[2].t3 106.907
R6782 ua[2].n23 ua[2].t9 106.907
R6783 ua[2].n0 ua[2].t0 87.3212
R6784 ua[2].n0 ua[2].t1 44.0792
R6785 ua[2].n27 ua[2] 4.89415
R6786 ua[2] ua[2].n26 2.98835
R6787 ua[2].n28 ua[2].n27 2.62026
R6788 ua[2].n27 ua[2] 2.53696
R6789 ua[2].n25 ua[2].n24 0.994487
R6790 ua[2].n26 ua[2].n25 0.592314
R6791 ua[2].n21 ua[2].n20 0.592314
R6792 ua[2].n17 ua[2].n16 0.592314
R6793 ua[2].n11 ua[2].n10 0.592314
R6794 ua[2].n9 ua[2].n8 0.592314
R6795 ua[2].n8 ua[2].n4 0.592314
R6796 ua[2].n12 ua[2].n11 0.592314
R6797 ua[2].n13 ua[2].n3 0.592314
R6798 ua[2].n14 ua[2].n13 0.592314
R6799 ua[2].n16 ua[2].n15 0.592314
R6800 ua[2].n19 ua[2].n18 0.592314
R6801 ua[2].n18 ua[2].n2 0.592314
R6802 ua[2].n22 ua[2].n21 0.592314
R6803 ua[2].n23 ua[2].n1 0.592314
R6804 ua[2].n24 ua[2].n23 0.592314
R6805 ua[2].n17 ua[2].n3 0.402674
R6806 ua[2].n15 ua[2].n14 0.402674
R6807 ua[2].n26 ua[2].n1 0.402674
R6808 ua[2].n10 ua[2].n9 0.394522
R6809 ua[2].n12 ua[2].n4 0.394522
R6810 ua[2].n6 ua[2].n4 0.389087
R6811 ua[2].n9 ua[2].n7 0.389087
R6812 ua[2].n20 ua[2].n19 0.389087
R6813 ua[2].n22 ua[2].n2 0.389087
R6814 ua[2].n24 ua[2].n22 0.378217
R6815 ua[2].n20 ua[2].n1 0.378217
R6816 ua[2].n14 ua[2].n12 0.372783
R6817 ua[2].n10 ua[2].n3 0.372783
R6818 ua[2].n7 ua[2].n5 0.36932
R6819 ua[2].n6 ua[2].n5 0.36932
R6820 ua[2].n15 ua[2].n2 0.356478
R6821 ua[2].n19 ua[2].n17 0.356478
R6822 ua[2] ua[2].n0 0.291805
R6823 ua[2].n28 ua[2] 0.0495889
R6824 ua[2] ua[2].n28 0.0493177
R6825 VCR_0.VT.n10 VCR_0.VT.t11 33.665
R6826 VCR_0.VT.n10 VCR_0.VT.t12 32.2761
R6827 VCR_0.VT.n4 VCR_0.VT.n3 17.3297
R6828 VCR_0.VT.n8 VCR_0.VT.n0 16.4338
R6829 VCR_0.VT.n7 VCR_0.VT.n1 16.4338
R6830 VCR_0.VT.n4 VCR_0.VT.n2 16.4338
R6831 VCR_0.VT.n6 VCR_0.VT.n5 16.4338
R6832 VCR_0.VT.n9 VCR_0.VT.t10 11.3457
R6833 VCR_0.VT.n0 VCR_0.VT.t6 3.3065
R6834 VCR_0.VT.n0 VCR_0.VT.t5 3.3065
R6835 VCR_0.VT.n1 VCR_0.VT.t4 3.3065
R6836 VCR_0.VT.n1 VCR_0.VT.t3 3.3065
R6837 VCR_0.VT.n2 VCR_0.VT.t8 3.3065
R6838 VCR_0.VT.n2 VCR_0.VT.t0 3.3065
R6839 VCR_0.VT.n3 VCR_0.VT.t2 3.3065
R6840 VCR_0.VT.n3 VCR_0.VT.t1 3.3065
R6841 VCR_0.VT.n5 VCR_0.VT.t7 3.3065
R6842 VCR_0.VT.n5 VCR_0.VT.t9 3.3065
R6843 VCR_0.VT VCR_0.VT.n10 1.23675
R6844 VCR_0.VT.n9 VCR_0.VT.n8 0.96925
R6845 VCR_0.VT.n8 VCR_0.VT.n7 0.896333
R6846 VCR_0.VT.n7 VCR_0.VT.n6 0.896333
R6847 VCR_0.VT.n6 VCR_0.VT.n4 0.896333
R6848 VCR_0.VT VCR_0.VT.n9 0.385917
R6849 a_6404_16954.n17 a_6404_16954.t1 25.6078
R6850 a_6404_16954.t0 a_6404_16954.n17 23.4966
R6851 a_6404_16954.n14 a_6404_16954.t3 23.2869
R6852 a_6404_16954.n7 a_6404_16954.t5 23.2869
R6853 a_6404_16954.n11 a_6404_16954.t7 15.6115
R6854 a_6404_16954.t7 a_6404_16954.n2 15.6115
R6855 a_6404_16954.n8 a_6404_16954.t4 15.6115
R6856 a_6404_16954.t4 a_6404_16954.n6 15.6115
R6857 a_6404_16954.n6 a_6404_16954.t6 15.6115
R6858 a_6404_16954.t6 a_6404_16954.n5 15.6115
R6859 a_6404_16954.n11 a_6404_16954.t2 15.6115
R6860 a_6404_16954.t2 a_6404_16954.n1 15.6115
R6861 a_6404_16954.n8 a_6404_16954.n2 8.48963
R6862 a_6404_16954.n5 a_6404_16954.n1 8.35104
R6863 a_6404_16954.n17 a_6404_16954.n16 7.9767
R6864 a_6404_16954.n8 a_6404_16954.n7 7.06613
R6865 a_6404_16954.n16 a_6404_16954.n0 6.56044
R6866 a_6404_16954.n5 a_6404_16954.n4 5.38843
R6867 a_6404_16954.n15 a_6404_16954.n1 4.29475
R6868 a_6404_16954.n4 a_6404_16954.t10 4.20487
R6869 a_6404_16954.n14 a_6404_16954.n13 3.72266
R6870 a_6404_16954.n3 a_6404_16954.t8 2.68574
R6871 a_6404_16954.n3 a_6404_16954.t9 2.68574
R6872 a_6404_16954.n11 a_6404_16954.n10 2.08746
R6873 a_6404_16954.n16 a_6404_16954.n15 1.77302
R6874 a_6404_16954.n7 a_6404_16954.n0 1.50128
R6875 a_6404_16954.n15 a_6404_16954.n14 1.50128
R6876 a_6404_16954.n6 a_6404_16954.n0 1.47643
R6877 a_6404_16954.n12 a_6404_16954.n1 0.223676
R6878 a_6404_16954.n10 a_6404_16954.n5 0.223676
R6879 a_6404_16954.n9 a_6404_16954.n8 0.223676
R6880 a_6404_16954.n13 a_6404_16954.n2 0.223676
R6881 a_6404_16954.n4 a_6404_16954.n3 0.116907
R6882 a_6404_16954.n9 a_6404_16954.n6 0.0455311
R6883 a_6404_16954.n12 a_6404_16954.n11 0.0300031
R6884 a_6404_16954.n10 a_6404_16954.n9 0.0136988
R6885 a_6404_16954.n13 a_6404_16954.n12 0.00709938
R6886 a_10404_14647.n2 a_10404_14647.t9 654.941
R6887 a_10404_14647.n2 a_10404_14647.t1 654.191
R6888 a_10404_14647.t0 a_10404_14647.n6 229.595
R6889 a_10404_14647.n0 a_10404_14647.t2 169.452
R6890 a_10404_14647.n0 a_10404_14647.t4 168.163
R6891 a_10404_14647.n1 a_10404_14647.t8 84.0197
R6892 a_10404_14647.n4 a_10404_14647.t6 23.2869
R6893 a_10404_14647.n4 a_10404_14647.t3 23.2869
R6894 a_10404_14647.n3 a_10404_14647.t7 23.2869
R6895 a_10404_14647.n3 a_10404_14647.t5 23.2869
R6896 a_10404_14647.n5 a_10404_14647.n2 7.85625
R6897 a_10404_14647.n6 a_10404_14647.n5 7.78276
R6898 a_10404_14647.n6 a_10404_14647.n1 6.26012
R6899 a_10404_14647.n1 a_10404_14647.n0 2.438
R6900 a_10404_14647.n4 a_10404_14647.n3 2.25174
R6901 a_10404_14647.n5 a_10404_14647.n4 1.04383
R6902 latch_sch_0.Qn.n1 latch_sch_0.Qn.t5 237.504
R6903 latch_sch_0.Qn.n3 latch_sch_0.Qn.t1 233.115
R6904 latch_sch_0.Qn.n1 latch_sch_0.Qn.t4 121.347
R6905 latch_sch_0.Qn.n0 latch_sch_0.Qn.t2 89.1813
R6906 latch_sch_0.Qn.n0 latch_sch_0.Qn.t3 87.4384
R6907 latch_sch_0.Qn.n2 latch_sch_0.Qn.n1 5.12424
R6908 latch_sch_0.Qn latch_sch_0.Qn.t0 4.88309
R6909 latch_sch_0.Qn.n2 latch_sch_0.Qn.n0 1.25771
R6910 latch_sch_0.Qn latch_sch_0.Qn.n3 0.516704
R6911 latch_sch_0.Qn.n3 latch_sch_0.Qn.n2 0.227352
R6912 a_21737_7899.t11 a_21737_7899.n13 301.625
R6913 a_21737_7899.n6 a_21737_7899.t4 301.625
R6914 a_21737_7899.n14 a_21737_7899.t11 300.925
R6915 a_21737_7899.t3 a_21737_7899.n1 300.925
R6916 a_21737_7899.n13 a_21737_7899.t3 300.925
R6917 a_21737_7899.t7 a_21737_7899.n11 300.925
R6918 a_21737_7899.n12 a_21737_7899.t7 300.925
R6919 a_21737_7899.n10 a_21737_7899.t8 300.925
R6920 a_21737_7899.t8 a_21737_7899.n2 300.925
R6921 a_21737_7899.n9 a_21737_7899.t5 300.925
R6922 a_21737_7899.t5 a_21737_7899.n8 300.925
R6923 a_21737_7899.t6 a_21737_7899.n3 300.925
R6924 a_21737_7899.n7 a_21737_7899.t6 300.925
R6925 a_21737_7899.t9 a_21737_7899.n5 300.925
R6926 a_21737_7899.n6 a_21737_7899.t9 300.925
R6927 a_21737_7899.n4 a_21737_7899.t4 300.925
R6928 a_21737_7899.n15 a_21737_7899.t1 96.0066
R6929 a_21737_7899.n0 a_21737_7899.t2 60.9515
R6930 a_21737_7899.n4 a_21737_7899.t10 23.0386
R6931 a_21737_7899.t0 a_21737_7899.n17 13.9376
R6932 a_21737_7899.n15 a_21737_7899.n0 1.80042
R6933 a_21737_7899.n16 a_21737_7899.n14 1.73148
R6934 a_21737_7899.n17 a_21737_7899.n16 0.996006
R6935 a_21737_7899.n13 a_21737_7899.n12 0.701587
R6936 a_21737_7899.n12 a_21737_7899.n2 0.701587
R6937 a_21737_7899.n8 a_21737_7899.n2 0.701587
R6938 a_21737_7899.n8 a_21737_7899.n7 0.701587
R6939 a_21737_7899.n7 a_21737_7899.n6 0.701587
R6940 a_21737_7899.n14 a_21737_7899.n1 0.701587
R6941 a_21737_7899.n11 a_21737_7899.n1 0.701587
R6942 a_21737_7899.n11 a_21737_7899.n10 0.701587
R6943 a_21737_7899.n10 a_21737_7899.n9 0.701587
R6944 a_21737_7899.n9 a_21737_7899.n3 0.701587
R6945 a_21737_7899.n5 a_21737_7899.n3 0.701587
R6946 a_21737_7899.n5 a_21737_7899.n4 0.611484
R6947 a_21737_7899.n16 a_21737_7899.n15 0.463884
R6948 a_21737_7899.n17 a_21737_7899.n0 0.248096
R6949 ua[0].n3 ua[0].n2 26.0898
R6950 ua[0].n6 ua[0].n5 25.7557
R6951 ua[0].n4 ua[0].n0 25.725
R6952 ua[0].n3 ua[0].n1 25.725
R6953 ua[0].n5 ua[0].t1 3.25874
R6954 ua[0].n5 ua[0].t6 3.25874
R6955 ua[0].n0 ua[0].t5 3.25874
R6956 ua[0].n0 ua[0].t4 3.25874
R6957 ua[0].n1 ua[0].t3 3.25874
R6958 ua[0].n1 ua[0].t2 3.25874
R6959 ua[0].n2 ua[0].t0 3.25874
R6960 ua[0].n2 ua[0].t7 3.25874
R6961 ua[0].n4 ua[0].n3 0.3755
R6962 ua[0].n6 ua[0].n4 0.345703
R6963 ua[0] ua[0].n6 0.301306
R6964 a_5453_6051.n0 a_5453_6051.t6 101.662
R6965 a_5453_6051.n0 a_5453_6051.t7 99.9341
R6966 a_5453_6051.t0 a_5453_6051.n12 91.9637
R6967 a_5453_6051.n1 a_5453_6051.t5 91.3528
R6968 a_5453_6051.n9 a_5453_6051.t4 82.8472
R6969 a_5453_6051.n4 a_5453_6051.t2 82.8472
R6970 a_5453_6051.n6 a_5453_6051.t8 49.4085
R6971 a_5453_6051.t10 a_5453_6051.n7 20.6938
R6972 a_5453_6051.n8 a_5453_6051.t10 20.6938
R6973 a_5453_6051.t9 a_5453_6051.n2 20.6938
R6974 a_5453_6051.n3 a_5453_6051.t9 20.6938
R6975 a_5453_6051.t3 a_5453_6051.n7 15.7488
R6976 a_5453_6051.t1 a_5453_6051.n2 15.7488
R6977 a_5453_6051.n8 a_5453_6051.t3 15.7488
R6978 a_5453_6051.n3 a_5453_6051.t1 15.7488
R6979 a_5453_6051.n6 a_5453_6051.n5 8.5685
R6980 a_5453_6051.n11 a_5453_6051.n10 7.9105
R6981 a_5453_6051.n1 a_5453_6051.n0 4.22661
R6982 a_5453_6051.n11 a_5453_6051.n6 2.39934
R6983 a_5453_6051.n9 a_5453_6051.n8 2.09913
R6984 a_5453_6051.n4 a_5453_6051.n3 2.09913
R6985 a_5453_6051.n12 a_5453_6051.n1 1.98693
R6986 a_5453_6051.n10 a_5453_6051.n7 1.90761
R6987 a_5453_6051.n5 a_5453_6051.n2 1.90761
R6988 a_5453_6051.n12 a_5453_6051.n11 0.160554
R6989 a_5453_6051.n10 a_5453_6051.n9 0.113336
R6990 a_5453_6051.n5 a_5453_6051.n4 0.113336
R6991 latch_sch_0.R.t3 latch_sch_0.R.t4 359.979
R6992 latch_sch_0.R latch_sch_0.R.t3 244.089
R6993 latch_sch_0.R.n0 latch_sch_0.R.t1 103.389
R6994 latch_sch_0.R.n0 latch_sch_0.R.t2 101.189
R6995 latch_sch_0.R.n1 latch_sch_0.R.t0 94.468
R6996 latch_sch_0.R.n1 latch_sch_0.R.n0 0.263273
R6997 latch_sch_0.R latch_sch_0.R.n1 0.163268
R6998 a_5453_6767.t0 a_5453_6767.n12 100.184
R6999 a_5453_6767.n12 a_5453_6767.t1 98.8091
R7000 a_5453_6767.n5 a_5453_6767.t3 97.2317
R7001 a_5453_6767.n5 a_5453_6767.t2 94.3099
R7002 a_5453_6767.n9 a_5453_6767.t5 82.8472
R7003 a_5453_6767.n2 a_5453_6767.t7 82.8472
R7004 a_5453_6767.n4 a_5453_6767.t10 51.083
R7005 a_5453_6767.t8 a_5453_6767.n7 20.6938
R7006 a_5453_6767.n8 a_5453_6767.t8 20.6938
R7007 a_5453_6767.t9 a_5453_6767.n0 20.6938
R7008 a_5453_6767.n1 a_5453_6767.t9 20.6938
R7009 a_5453_6767.t4 a_5453_6767.n7 15.7488
R7010 a_5453_6767.t6 a_5453_6767.n0 15.7488
R7011 a_5453_6767.n8 a_5453_6767.t4 15.7488
R7012 a_5453_6767.n1 a_5453_6767.t6 15.7488
R7013 a_5453_6767.n4 a_5453_6767.n3 11.9173
R7014 a_5453_6767.n11 a_5453_6767.n10 11.8323
R7015 a_5453_6767.n12 a_5453_6767.n11 3.79321
R7016 a_5453_6767.n11 a_5453_6767.n6 2.28765
R7017 a_5453_6767.n2 a_5453_6767.n1 2.09913
R7018 a_5453_6767.n9 a_5453_6767.n8 2.09848
R7019 a_5453_6767.n10 a_5453_6767.n7 1.92106
R7020 a_5453_6767.n3 a_5453_6767.n0 1.90761
R7021 a_5453_6767.n6 a_5453_6767.n4 0.464091
R7022 a_5453_6767.n6 a_5453_6767.n5 0.175682
R7023 a_5453_6767.n10 a_5453_6767.n9 0.113336
R7024 a_5453_6767.n3 a_5453_6767.n2 0.113336
R7025 a_20802_14722.t0 a_20802_14722.n1 657.601
R7026 a_20802_14722.n1 a_20802_14722.n0 4.96288
R7027 a_20802_14722.n1 a_20802_14722.t2 4.03765
R7028 a_20802_14722.n0 a_20802_14722.t1 0.0629965
R7029 a_20802_14722.n0 a_20802_14722.t3 0.0586811
R7030 COMP_2_0.vin_n.n0 COMP_2_0.vin_n.t0 233.142
R7031 COMP_2_0.vin_n.n0 COMP_2_0.vin_n.t1 231.877
R7032 COMP_2_0.vin_n.n1 COMP_2_0.vin_n.t2 33.601
R7033 COMP_2_0.vin_n.n1 COMP_2_0.vin_n.t3 32.2522
R7034 COMP_2_0.vin_n COMP_2_0.vin_n.n0 3.77777
R7035 COMP_2_0.vin_n COMP_2_0.vin_n.n1 0.771552
R7036 a_6061_11160.n0 a_6061_11160.t4 118.172
R7037 a_6061_11160.t1 a_6061_11160.n1 96.5512
R7038 a_6061_11160.n0 a_6061_11160.t3 96.5491
R7039 a_6061_11160.n0 a_6061_11160.t0 96.5469
R7040 a_6061_11160.n1 a_6061_11160.t2 96.5448
R7041 a_6061_11160.n1 a_6061_11160.n0 0.663044
R7042 delay_1_0.vd_n.n3 delay_1_0.vd_n.t0 238.923
R7043 delay_1_0.vd_n delay_1_0.vd_n.n4 18.3251
R7044 delay_1_0.vd_n.n4 delay_1_0.vd_n 7.08575
R7045 delay_1_0.vd_n delay_1_0.vd_n.t1 6.86073
R7046 delay_1_0.vd_n delay_1_0.vd_n.t5 6.68369
R7047 delay_1_0.vd_n.n4 delay_1_0.vd_n 5.26786
R7048 delay_1_0.vd_n delay_1_0.vd_n.n3 0.259595
R7049 delay_1_0.vd_n.n2 delay_1_0.vd_n.n1 0.215474
R7050 delay_1_0.vd_n.n3 delay_1_0.vd_n.n2 0.136892
R7051 delay_1_0.vd_n.n1 delay_1_0.vd_n.t3 0.092145
R7052 delay_1_0.vd_n.n0 delay_1_0.vd_n.t6 0.0918192
R7053 delay_1_0.vd_n.n2 delay_1_0.vd_n.n0 0.0197857
R7054 delay_1_0.vd_n.n1 delay_1_0.vd_n.t2 0.00132177
R7055 delay_1_0.vd_n.n0 delay_1_0.vd_n.t4 0.00132177
R7056 ua[3] ua[3].n0 9.21498
R7057 ua[3].n0 ua[3].t2 4.66216
R7058 ua[3].n0 ua[3].t0 4.66216
R7059 ua[3].n0 ua[3].t1 4.66216
R7060 a_11329_22619.t0 a_11329_22619.n12 668.698
R7061 a_11329_22619.n10 a_11329_22619.t1 31.4954
R7062 a_11329_22619.n9 a_11329_22619.t6 30.0086
R7063 a_11329_22619.n3 a_11329_22619.t4 29.798
R7064 a_11329_22619.n10 a_11329_22619.t2 26.5479
R7065 a_11329_22619.n11 a_11329_22619.n10 9.04454
R7066 a_11329_22619.n6 a_11329_22619.t7 8.67282
R7067 a_11329_22619.n1 a_11329_22619.t8 8.34339
R7068 a_11329_22619.n4 a_11329_22619.n3 5.50673
R7069 a_11329_22619.n12 a_11329_22619.n11 4.918
R7070 a_11329_22619.n5 a_11329_22619.n4 3.96009
R7071 a_11329_22619.n8 a_11329_22619.n7 3.62746
R7072 a_11329_22619.n4 a_11329_22619.t3 3.59247
R7073 a_11329_22619.n8 a_11329_22619.t5 3.53527
R7074 a_11329_22619.n11 a_11329_22619.n9 2.90932
R7075 a_11329_22619.n9 a_11329_22619.n8 2.54528
R7076 a_11329_22619.n12 a_11329_22619.n0 2.36329
R7077 a_11329_22619.n7 a_11329_22619.n6 0.53261
R7078 a_11329_22619.n2 a_11329_22619.n1 0.494766
R7079 a_11329_22619.n3 a_11329_22619.n0 0.413242
R7080 a_11329_22619.n2 a_11329_22619.n0 0.324367
R7081 a_11329_22619.n7 a_11329_22619.n1 0.312375
R7082 a_11329_22619.n6 a_11329_22619.n5 0.312375
R7083 a_11329_22619.n5 a_11329_22619.n2 0.038344
R7084 COMP_2_0.vb.n6 COMP_2_0.vb.t3 227.369
R7085 COMP_2_0.vb.n7 COMP_2_0.vb.t0 169.452
R7086 COMP_2_0.vb.n7 COMP_2_0.vb.t1 168.163
R7087 COMP_2_0.vb.n8 COMP_2_0.vb.n6 8.71954
R7088 COMP_2_0.vb COMP_2_0.vb.t9 6.22797
R7089 COMP_2_0.vb.n0 COMP_2_0.vb.t10 5.60946
R7090 COMP_2_0.vb.n3 COMP_2_0.vb.t4 3.56652
R7091 COMP_2_0.vb.n5 COMP_2_0.vb.n4 3.54337
R7092 COMP_2_0.vb.n4 COMP_2_0.vb.t5 3.0689
R7093 COMP_2_0.vb.n2 COMP_2_0.vb.n1 2.86516
R7094 COMP_2_0.vb.n4 COMP_2_0.vb.n3 2.85956
R7095 COMP_2_0.vb.n1 COMP_2_0.vb.n0 2.85912
R7096 COMP_2_0.vb.n3 COMP_2_0.vb.n2 2.85912
R7097 COMP_2_0.vb.n0 COMP_2_0.vb.t8 2.69352
R7098 COMP_2_0.vb.n2 COMP_2_0.vb.t7 2.69352
R7099 COMP_2_0.vb.n1 COMP_2_0.vb.t6 2.69273
R7100 COMP_2_0.vb.n5 COMP_2_0.vb.t2 2.02902
R7101 COMP_2_0.vb.n6 COMP_2_0.vb.n5 1.36824
R7102 COMP_2_0.vb.n8 COMP_2_0.vb.n7 1.22406
R7103 COMP_2_0.vb COMP_2_0.vb.n8 1.05098
R7104 ua[4].t1 ua[4].t2 18.6605
R7105 ua[4].t0 ua[4].t1 18.6605
R7106 ua[4] ua[4].t0 13.672
R7107 BIAS_1_0.XQ4.Emitter.n17 BIAS_1_0.XQ4.Emitter.n12 83.5719
R7108 BIAS_1_0.XQ4.Emitter.n16 BIAS_1_0.XQ4.Emitter.n14 83.5719
R7109 BIAS_1_0.XQ4.Emitter.n15 BIAS_1_0.XQ4.Emitter.n0 83.5719
R7110 BIAS_1_0.XQ4.Emitter.n15 BIAS_1_0.XQ4.Emitter.n4 73.3165
R7111 BIAS_1_0.XQ4.Emitter.n18 BIAS_1_0.XQ4.Emitter.n17 73.19
R7112 BIAS_1_0.XQ4.Emitter.n1 BIAS_1_0.XQ4.Emitter.t1 38.8946
R7113 BIAS_1_0.XQ4.Emitter.n1 BIAS_1_0.XQ4.Emitter.t0 31.7107
R7114 BIAS_1_0.XQ4.Emitter.n16 BIAS_1_0.XQ4.Emitter.n15 26.074
R7115 BIAS_1_0.XQ4.Emitter.n17 BIAS_1_0.XQ4.Emitter.t2 25.7843
R7116 BIAS_1_0.XQ4.Emitter.n13 BIAS_1_0.XQ4.Emitter.n8 9.3005
R7117 BIAS_1_0.XQ4.Emitter.n23 BIAS_1_0.XQ4.Emitter.n13 9.3005
R7118 BIAS_1_0.XQ4.Emitter.n13 BIAS_1_0.XQ4.Emitter.n9 9.3005
R7119 BIAS_1_0.XQ4.Emitter.n13 BIAS_1_0.XQ4.Emitter.n10 9.3005
R7120 BIAS_1_0.XQ4.Emitter.n22 BIAS_1_0.XQ4.Emitter.n8 9.3005
R7121 BIAS_1_0.XQ4.Emitter.n23 BIAS_1_0.XQ4.Emitter.n22 9.3005
R7122 BIAS_1_0.XQ4.Emitter.n22 BIAS_1_0.XQ4.Emitter.n9 9.3005
R7123 BIAS_1_0.XQ4.Emitter.n22 BIAS_1_0.XQ4.Emitter.n10 9.3005
R7124 BIAS_1_0.XQ4.Emitter.n10 BIAS_1_0.XQ4.Emitter.n3 9.3005
R7125 BIAS_1_0.XQ4.Emitter.n25 BIAS_1_0.XQ4.Emitter.n3 9.3005
R7126 BIAS_1_0.XQ4.Emitter.n9 BIAS_1_0.XQ4.Emitter.n3 9.3005
R7127 BIAS_1_0.XQ4.Emitter.n23 BIAS_1_0.XQ4.Emitter.n3 9.3005
R7128 BIAS_1_0.XQ4.Emitter.n10 BIAS_1_0.XQ4.Emitter.n6 9.3005
R7129 BIAS_1_0.XQ4.Emitter.n25 BIAS_1_0.XQ4.Emitter.n6 9.3005
R7130 BIAS_1_0.XQ4.Emitter.n9 BIAS_1_0.XQ4.Emitter.n6 9.3005
R7131 BIAS_1_0.XQ4.Emitter.n23 BIAS_1_0.XQ4.Emitter.n6 9.3005
R7132 BIAS_1_0.XQ4.Emitter.n10 BIAS_1_0.XQ4.Emitter.n2 9.3005
R7133 BIAS_1_0.XQ4.Emitter.n25 BIAS_1_0.XQ4.Emitter.n2 9.3005
R7134 BIAS_1_0.XQ4.Emitter.n9 BIAS_1_0.XQ4.Emitter.n2 9.3005
R7135 BIAS_1_0.XQ4.Emitter.n23 BIAS_1_0.XQ4.Emitter.n2 9.3005
R7136 BIAS_1_0.XQ4.Emitter.n8 BIAS_1_0.XQ4.Emitter.n2 9.3005
R7137 BIAS_1_0.XQ4.Emitter.n24 BIAS_1_0.XQ4.Emitter.n10 9.3005
R7138 BIAS_1_0.XQ4.Emitter.n25 BIAS_1_0.XQ4.Emitter.n24 9.3005
R7139 BIAS_1_0.XQ4.Emitter.n24 BIAS_1_0.XQ4.Emitter.n9 9.3005
R7140 BIAS_1_0.XQ4.Emitter.n24 BIAS_1_0.XQ4.Emitter.n8 9.3005
R7141 BIAS_1_0.XQ4.Emitter.n24 BIAS_1_0.XQ4.Emitter.n23 9.3005
R7142 BIAS_1_0.XQ4.Emitter.n2 BIAS_1_0.XQ4.Emitter.n1 4.95643
R7143 BIAS_1_0.XQ4.Emitter.n25 BIAS_1_0.XQ4.Emitter.n5 4.64588
R7144 BIAS_1_0.XQ4.Emitter.n21 BIAS_1_0.XQ4.Emitter.n20 4.64588
R7145 BIAS_1_0.XQ4.Emitter.n8 BIAS_1_0.XQ4.Emitter.n7 4.64588
R7146 BIAS_1_0.XQ4.Emitter.n20 BIAS_1_0.XQ4.Emitter.n19 4.64588
R7147 BIAS_1_0.XQ4.Emitter.n20 BIAS_1_0.XQ4.Emitter.n11 4.64588
R7148 BIAS_1_0.XQ4.Emitter.n12 BIAS_1_0.XQ4.Emitter.n8 1.25468
R7149 BIAS_1_0.XQ4.Emitter.n25 BIAS_1_0.XQ4.Emitter.n4 1.19225
R7150 BIAS_1_0.XQ4.Emitter.n23 BIAS_1_0.XQ4.Emitter.n14 1.07024
R7151 BIAS_1_0.XQ4.Emitter.n18 BIAS_1_0.XQ4.Emitter.n8 1.0237
R7152 BIAS_1_0.XQ4.Emitter.n9 BIAS_1_0.XQ4.Emitter.n0 0.885803
R7153 BIAS_1_0.XQ4.Emitter.n20 BIAS_1_0.XQ4.Emitter.n18 0.812055
R7154 BIAS_1_0.XQ4.Emitter.n14 BIAS_1_0.XQ4.Emitter.n9 0.77514
R7155 BIAS_1_0.XQ4.Emitter BIAS_1_0.XQ4.Emitter.n0 0.756696
R7156 BIAS_1_0.XQ4.Emitter.n10 BIAS_1_0.XQ4.Emitter.n4 0.647417
R7157 BIAS_1_0.XQ4.Emitter.n23 BIAS_1_0.XQ4.Emitter.n12 0.590702
R7158 BIAS_1_0.XQ4.Emitter.t2 BIAS_1_0.XQ4.Emitter.n16 0.290206
R7159 BIAS_1_0.XQ4.Emitter BIAS_1_0.XQ4.Emitter.n25 0.203382
R7160 BIAS_1_0.XQ4.Emitter.n24 BIAS_1_0.XQ4.Emitter.n11 0.0112346
R7161 BIAS_1_0.XQ4.Emitter.n22 BIAS_1_0.XQ4.Emitter.n5 0.0112346
R7162 BIAS_1_0.XQ4.Emitter.n21 BIAS_1_0.XQ4.Emitter.n3 0.0112346
R7163 BIAS_1_0.XQ4.Emitter.n7 BIAS_1_0.XQ4.Emitter.n6 0.0112346
R7164 BIAS_1_0.XQ4.Emitter.n19 BIAS_1_0.XQ4.Emitter.n2 0.0112346
R7165 BIAS_1_0.XQ4.Emitter.n13 BIAS_1_0.XQ4.Emitter.n11 0.0112346
R7166 BIAS_1_0.XQ4.Emitter.n13 BIAS_1_0.XQ4.Emitter.n5 0.0112346
R7167 BIAS_1_0.XQ4.Emitter.n22 BIAS_1_0.XQ4.Emitter.n21 0.0112346
R7168 BIAS_1_0.XQ4.Emitter.n7 BIAS_1_0.XQ4.Emitter.n3 0.0112346
R7169 BIAS_1_0.XQ4.Emitter.n19 BIAS_1_0.XQ4.Emitter.n6 0.0112346
R7170 ua[1].n3 ua[1].t1 34.4698
R7171 ua[1].t1 ua[1].n1 34.4692
R7172 ua[1].n2 ua[1].t0 17.1948
R7173 ua[1].n2 ua[1].n0 3.01859
R7174 ua[1].n5 ua[1].n0 2.41294
R7175 ua[1].n3 ua[1].n2 1.40867
R7176 ua[1].n1 ua[1].n0 0.9005
R7177 ua[1] ua[1].n5 0.67231
R7178 ua[1].n5 ua[1].n4 0.301078
R7179 ua[1].n4 ua[1].n3 0.166107
R7180 ua[1].n4 ua[1].n1 0.00100004
C0 a_17267_7131# a_15577_6765# 0
C1 a_14689_10265# a_14097_10265# 0.06616f
C2 a_9886_27451# a_9886_27747# 0.16485f
C3 a_17853_5073# a_17267_4669# 0.0513f
C4 latch_sch_0.Qn latch_sch_0.R 0.35822f
C5 latch_sch_0.R a_12495_10665# 0.1132f
C6 a_9886_27747# delay_1_0.vd_n 0
C7 a_4266_30348# a_3674_30348# 0.06471f
C8 ua[2] ua[4] 0.2849f
C9 latch_sch_0.Qn a_3674_30348# 0.00395f
C10 a_6064_20056# COMP_2_0.vb 0.75714f
C11 a_16681_5073# ua[4] 0.01487f
C12 a_11336_20947# VAPWR 0
C13 a_14985_6107# a_15577_6107# 0.06621f
C14 a_14985_6765# a_14393_6765# 0.06623f
C15 a_14985_6765# ua[3] 0
C16 ua[2] a_19010_2607# 0.10565f
C17 a_9886_25971# a_9886_26267# 0.16485f
C18 a_12844_27155# a_12844_26563# 0.06471f
C19 a_14097_6107# a_14393_6765# 0.06573f
C20 COMP_2_0.vin_n VCR_0.VT 1.90539f
C21 BIAS_1_0.XQ12.Emitter delay_1_0.vd_n 0.00471f
C22 delay_1_0.vd_n COMP_2_0.vb 0.53503f
C23 ua[1] VAPWR 0.05767f
C24 latch_sch_0.Qn Timming_0.Vd 0.98025f
C25 Timming_0.Vd a_12495_10665# 0.03805f
C26 a_17267_7131# Timming_0.Vd 0
C27 a_17853_5073# ua[4] 0.06831f
C28 a_14985_6765# a_15577_6765# 0.06625f
C29 ua[0] a_21737_3791# 0.00365f
C30 a_15281_10265# a_14689_10265# 0.06624f
C31 a_4858_30348# a_5450_30348# 0.06668f
C32 a_8096_19998# a_9068_19998# 0.00723f
C33 a_11336_20947# BIAS_1_0.XQ4.Emitter 0.29657f
C34 a_7124_24056# COMP_2_0.vb 0.25529f
C35 ua[5] ua[4] 0.03264f
C36 a_12844_27155# BIAS_1_0.XQ12.Emitter 0.07519f
C37 a_17853_5073# a_19010_2607# 0.129f
C38 a_5154_35748# a_4858_35748# 0.16485f
C39 ua[4] VCR_0.VT 0.11395f
C40 a_2786_41806# a_3378_41806# 0.06471f
C41 ua[2] a_21737_3791# 0.0014f
C42 a_9554_24056# COMP_2_0.vb 0.2233f
C43 latch_sch_0.Qn a_12179_10665# 0.03721f
C44 VAPWR latch_sch_0.R 2.14354f
C45 latch_sch_0.Qn COMP_2_0.vb 0.1384f
C46 a_15577_6765# ua[3] 0.00218f
C47 a_9886_27451# a_9886_27155# 0.16485f
C48 a_18714_5807# ua[3] 0.03238f
C49 a_16169_6107# ua[3] 0.10237f
C50 a_14985_6765# Timming_0.Vd 0.00295f
C51 a_3082_35748# a_3378_35748# 0.16485f
C52 ua[2] a_16681_2611# 0.0165f
C53 VAPWR a_8279_30718# 0.25761f
C54 a_11336_20947# a_12844_26563# 0
C55 VAPWR Timming_0.Vd 1.34646f
C56 a_4266_30348# a_4858_30348# 0.06471f
C57 latch_sch_0.Qn ua[5] 0.59877f
C58 ua[0] VAPWR 6.15268f
C59 a_9886_25379# COMP_2_0.vb 0
C60 a_14689_2607# a_14097_2607# 0.06619f
C61 a_14393_6107# a_14985_6107# 0.06618f
C62 a_14393_6765# Timming_0.Vd 0
C63 ua[3] Timming_0.Vd 0.05857f
C64 ua[1] ua[0] 0
C65 a_17267_4669# ua[4] 0.25912f
C66 a_7586_25675# a_7586_26267# 0.06471f
C67 COMP_2_0.vin_n a_6064_20056# 0.28782f
C68 a_11336_20947# BIAS_1_0.XQ12.Emitter 0.01756f
C69 a_11336_20947# COMP_2_0.vb 0.32832f
C70 a_19306_5807# ua[3] 0.00102f
C71 VAPWR a_12179_10665# 0.07679f
C72 a_15577_6765# Timming_0.Vd 0.09155f
C73 ua[2] ua[1] 0.25655f
C74 VAPWR COMP_2_0.vb 12.3003f
C75 COMP_2_0.vin_n delay_1_0.vd_n 0.58484f
C76 a_11336_20947# a_12844_25971# 0.0012f
C77 ua[2] ua[3] 0.26213f
C78 a_16169_6107# Timming_0.Vd 0.02545f
C79 ua[1] a_21737_5649# 1.90949f
C80 a_15577_6107# ua[3] 0.00215f
C81 latch_sch_0.R Timming_0.Vd 0.40879f
C82 a_16681_5073# ua[3] 0.37832f
C83 COMP_2_0.vb a_8582_24056# 0.22294f
C84 a_16681_2611# VCR_0.VT 0
C85 COMP_2_0.vin_n a_7124_24056# 0.0068f
C86 VAPWR a_10040_19998# 0.00872f
C87 a_18714_5807# a_19306_5807# 0.06742f
C88 latch_sch_0.Qn a_3082_30348# 0.08528f
C89 a_5450_30348# delay_1_0.vd_n 0.0073f
C90 a_3970_35748# a_4266_35748# 0.16485f
C91 a_15577_6107# a_15577_6765# 0.05493f
C92 BIAS_1_0.XQ12.Emitter BIAS_1_0.XQ4.Emitter 0.34399f
C93 a_19010_2607# ua[4] 0.00115f
C94 a_6064_20056# delay_1_0.vd_n 0.02898f
C95 ua[1] a_17853_5073# 0.03559f
C96 VAPWR ua[5] 0.52413f
C97 a_3970_41806# a_3378_41806# 0.06471f
C98 a_17853_5073# ua[3] 0.24362f
C99 a_9886_25379# a_9886_25675# 0.16485f
C100 a_16169_6107# a_15577_6107# 0.07401f
C101 COMP_2_0.vin_n latch_sch_0.Qn 0.1665f
C102 a_16169_6107# a_16681_5073# 0.05421f
C103 VAPWR a_4858_30348# 0
C104 a_9886_25971# a_9886_25675# 0.16485f
C105 latch_sch_0.R COMP_2_0.vb 0.03217f
C106 VAPWR VCR_0.VT 3.23544f
C107 a_15281_2607# ua[4] 0.001f
C108 a_6064_20056# a_7124_24056# 0.06762f
C109 a_5154_35748# a_5450_35748# 0.16485f
C110 a_9886_25379# a_9886_25083# 0.16485f
C111 ua[1] VCR_0.VT 0.26427f
C112 a_4266_30348# a_5450_30348# 0
C113 ua[3] VCR_0.VT 0.0586f
C114 a_7586_26859# a_7586_27451# 0.06471f
C115 a_17853_5073# a_18714_5807# 0.0126f
C116 latch_sch_0.R a_14097_10265# 0
C117 a_15873_10265# Timming_0.Vd 0.00258f
C118 a_7586_25675# a_7586_25083# 0.06471f
C119 Timming_0.Vd a_12179_10665# 0.11917f
C120 VAPWR a_8096_19998# 0.00557f
C121 a_9886_26563# a_9886_26267# 0.16485f
C122 BIAS_1_0.XQ12.Emitter a_12844_26563# 0.00162f
C123 a_14393_6107# a_14097_6107# 0.06576f
C124 ua[5] latch_sch_0.R 0.1913f
C125 a_11336_20947# a_12844_25379# 0.07245f
C126 a_6638_19998# COMP_2_0.vb 0.05342f
C127 latch_sch_0.Qn delay_1_0.vd_n 0.26098f
C128 a_12844_25971# a_12844_26563# 0.06471f
C129 latch_sch_0.R VCR_0.VT 0
C130 a_4266_35748# a_4562_35748# 0.16485f
C131 VAPWR a_9068_19998# 0.00548f
C132 a_9886_27155# a_9886_26859# 0.16485f
C133 a_15873_2607# ua[4] 0.04362f
C134 a_16681_2611# ua[4] 0.25834f
C135 COMP_2_0.vin_n VAPWR 3.09341f
C136 a_14393_6107# a_14393_6765# 0.05493f
C137 a_9886_26859# a_9886_26563# 0.16485f
C138 ua[5] Timming_0.Vd 0.41709f
C139 a_17267_4669# ua[3] 0.02205f
C140 a_3970_35748# a_3674_35748# 0.16485f
C141 a_17853_5073# a_19306_5807# 0.01401f
C142 BIAS_1_0.XQ12.Emitter a_12844_25971# 0
C143 latch_sch_0.Qn a_4266_30348# 0
C144 a_14985_6107# a_14985_6765# 0.05493f
C145 a_2786_35748# a_3082_35748# 0.16485f
C146 ua[2] a_17853_5073# 0.06751f
C147 VAPWR a_5450_30348# 0.42558f
C148 a_10040_19998# COMP_2_0.vb 0.13513f
C149 ua[0] VCR_0.VT 0.00365f
C150 latch_sch_0.Qn a_12495_10665# 0.11687f
C151 a_15281_2607# a_15873_2607# 0.06618f
C152 a_16681_2611# a_15281_2607# 0
C153 a_16169_6107# a_14393_6107# 0
C154 a_16681_5073# a_17853_5073# 0.02151f
C155 a_6064_20056# VAPWR 0.68144f
C156 a_3082_30348# a_3674_30348# 0.06471f
C157 a_16169_6107# a_17267_4669# 0.01369f
C158 ua[5] a_12179_10665# 0.11434f
C159 a_7586_26859# a_7586_26267# 0.06471f
C160 a_4562_41806# a_5154_41806# 0.06471f
C161 ua[2] VCR_0.VT 6.89088f
C162 ua[3] ua[4] 1.12519f
C163 VAPWR delay_1_0.vd_n 15.6496f
C164 a_14985_6107# ua[3] 0
C165 VCR_0.VT COMP_2_0.vb 0.01459f
C166 a_4562_35748# a_4858_35748# 0.16485f
C167 a_15281_10265# a_15873_10265# 0.06625f
C168 a_16169_6107# ua[4] 0.08219f
C169 a_5450_30348# a_3674_30348# 0
C170 a_17853_5073# VCR_0.VT 0
C171 COMP_2_0.vb a_8096_19998# 0.14251f
C172 a_7124_24056# a_8582_24056# 0.00723f
C173 a_16681_2611# a_15873_2607# 0.00527f
C174 a_16169_6107# a_14985_6107# 0
C175 VAPWR a_4266_30348# 0
C176 ua[5] VCR_0.VT 1.04093f
C177 latch_sch_0.Qn VAPWR 2.12045f
C178 VAPWR a_12495_10665# 0.07786f
C179 a_9886_25083# COMP_2_0.vb 0
C180 a_14689_2607# ua[4] 0
C181 a_3970_41806# a_4562_41806# 0.06471f
C182 a_9554_24056# a_8582_24056# 0.00723f
C183 a_3378_35748# a_3674_35748# 0.16485f
C184 ua[1] a_21737_3791# 0.84893f
C185 a_16681_5073# a_17267_4669# 0.04951f
C186 a_17267_7131# ua[3] 0.38354f
C187 COMP_2_0.vb a_9068_19998# 0.13517f
C188 a_7586_27451# delay_1_0.vd_n 0
C189 COMP_2_0.vin_n COMP_2_0.vb 0.93534f
C190 a_12844_25971# a_12844_25379# 0.06471f
C191 a_6064_20056# a_6638_19998# 0.14296f
C192 a_14689_2607# a_15281_2607# 0.06623f
C193 a_10040_19998# a_9068_19998# 0.00723f
C194 a_7586_25083# COMP_2_0.vb 0
C195 ua[0] VGND 7.21026f
C196 ua[1] VGND 19.3533f
C197 ua[2] VGND 20.32121f
C198 ua[4] VGND 19.1473f
C199 ua[3] VGND 18.7448f
C200 ua[5] VGND 7.34895f
C201 VAPWR VGND 0.35588p
C202 a_21737_3791# VGND 4.13855f
C203 a_21737_5649# VGND 4.40137f
C204 a_19306_5807# VGND 1.25829f
C205 a_19010_2607# VGND 1.20194f
C206 a_18714_5807# VGND 1.21224f
C207 a_17267_4669# VGND 0.47073f
C208 a_16681_2611# VGND 0.70042f
C209 a_17853_5073# VGND 2.70189f
C210 a_17267_7131# VGND 0.58358f
C211 a_16681_5073# VGND 0.41501f
C212 a_16169_6107# VGND 1.64417f
C213 a_15873_2607# VGND 1.24818f
C214 a_15577_6107# VGND 1.07044f
C215 a_15281_2607# VGND 1.23243f
C216 a_14985_6107# VGND 1.0715f
C217 a_14689_2607# VGND 1.23243f
C218 a_14393_6107# VGND 1.07199f
C219 a_14097_2607# VGND 1.31315f
C220 a_15873_10265# VGND 1.24245f
C221 a_15577_6765# VGND 1.07214f
C222 a_15281_10265# VGND 1.17504f
C223 a_14985_6765# VGND 1.07156f
C224 a_14689_10265# VGND 1.17504f
C225 a_14393_6765# VGND 1.07206f
C226 a_14097_6107# VGND 1.25481f
C227 a_14097_10265# VGND 1.25536f
C228 a_12495_10665# VGND 0.01639f
C229 a_12179_10665# VGND 0.01513f
C230 Timming_0.Vd VGND 19.26188f
C231 latch_sch_0.R VGND 4.81582f
C232 VCR_0.VT VGND 26.44499f
C233 a_10040_19998# VGND 0.61197f
C234 a_9554_24056# VGND 0.61994f
C235 a_9068_19998# VGND 0.60213f
C236 a_8582_24056# VGND 0.61279f
C237 a_8096_19998# VGND 0.61344f
C238 COMP_2_0.vb VGND 89.46873f
C239 a_7124_24056# VGND 1.09689f
C240 a_6638_19998# VGND 0.58617f
C241 a_6064_20056# VGND 35.9904f
C242 COMP_2_0.vin_n VGND 9.23523f
C243 a_11336_20947# VGND 9.36805f
C244 a_9886_25083# VGND 1.40376f
C245 a_9886_25379# VGND 1.28117f
C246 a_7586_25083# VGND 1.42009f
C247 BIAS_1_0.XQ4.Emitter VGND 5.7438f
C248 a_12844_25379# VGND 1.37614f
C249 a_9886_25675# VGND 1.31211f
C250 a_9886_25971# VGND 1.23556f
C251 a_7586_25675# VGND 1.36794f
C252 a_12844_25971# VGND 1.3281f
C253 a_9886_26267# VGND 1.25409f
C254 a_9886_26563# VGND 1.27876f
C255 a_7586_26267# VGND 1.36088f
C256 a_12844_26563# VGND 1.36088f
C257 a_9886_26859# VGND 1.27902f
C258 a_9886_27155# VGND 1.28083f
C259 a_7586_26859# VGND 1.37376f
C260 a_12844_27155# VGND 1.36228f
C261 a_9886_27451# VGND 1.27983f
C262 BIAS_1_0.XQ12.Emitter VGND 15.4118f
C263 a_9886_27747# VGND 1.45229f
C264 a_7586_27451# VGND 1.45159f
C265 delay_1_0.vd_n VGND 0.34507p
C266 a_8279_30718# VGND 0.35164f
C267 a_5450_30348# VGND 1.30048f
C268 a_4858_30348# VGND 1.18378f
C269 a_4266_30348# VGND 1.18164f
C270 a_3674_30348# VGND 1.18277f
C271 a_3082_30348# VGND 1.18319f
C272 latch_sch_0.Qn VGND 17.6584f
C273 a_5450_35748# VGND 1.36439f
C274 a_5154_35748# VGND 1.01786f
C275 a_5154_41806# VGND 1.30144f
C276 a_4858_35748# VGND 1.01781f
C277 a_4562_35748# VGND 1.0178f
C278 a_4562_41806# VGND 1.16107f
C279 a_4266_35748# VGND 1.0178f
C280 a_3970_35748# VGND 1.0178f
C281 a_3970_41806# VGND 1.16105f
C282 a_3674_35748# VGND 1.0178f
C283 a_3378_35748# VGND 1.01781f
C284 a_3378_41806# VGND 1.16107f
C285 a_3082_35748# VGND 1.01785f
C286 a_2786_35748# VGND 1.34385f
C287 a_2786_41806# VGND 1.29323f
C288 BIAS_1_0.XQ4.Emitter.n0 VGND 0.03776f
C289 BIAS_1_0.XQ4.Emitter.t1 VGND 0.12205f
C290 BIAS_1_0.XQ4.Emitter.t0 VGND 0.04158f
C291 BIAS_1_0.XQ4.Emitter.n1 VGND 0.94859f
C292 BIAS_1_0.XQ4.Emitter.n2 VGND 0.36198f
C293 BIAS_1_0.XQ4.Emitter.n3 VGND 0.07459f
C294 BIAS_1_0.XQ4.Emitter.n4 VGND 0.07743f
C295 BIAS_1_0.XQ4.Emitter.n6 VGND 0.07459f
C296 BIAS_1_0.XQ4.Emitter.n8 VGND 0.06379f
C297 BIAS_1_0.XQ4.Emitter.n9 VGND 0.03819f
C298 BIAS_1_0.XQ4.Emitter.n10 VGND 0.13664f
C299 BIAS_1_0.XQ4.Emitter.n12 VGND 0.04243f
C300 BIAS_1_0.XQ4.Emitter.n13 VGND 0.07459f
C301 BIAS_1_0.XQ4.Emitter.n14 VGND 0.04243f
C302 BIAS_1_0.XQ4.Emitter.n15 VGND 0.16991f
C303 BIAS_1_0.XQ4.Emitter.n16 VGND 0.03783f
C304 BIAS_1_0.XQ4.Emitter.t2 VGND 0.03742f
C305 BIAS_1_0.XQ4.Emitter.n17 VGND 0.17004f
C306 BIAS_1_0.XQ4.Emitter.n18 VGND 0.06974f
C307 BIAS_1_0.XQ4.Emitter.n20 VGND 0.13222f
C308 BIAS_1_0.XQ4.Emitter.n22 VGND 0.07459f
C309 BIAS_1_0.XQ4.Emitter.n23 VGND 0.03819f
C310 BIAS_1_0.XQ4.Emitter.n24 VGND 0.0731f
C311 BIAS_1_0.XQ4.Emitter.n25 VGND 0.03827f
C312 COMP_2_0.vb.t3 VGND 0.00297f
C313 COMP_2_0.vb.t5 VGND 0.71042f
C314 COMP_2_0.vb.t4 VGND 0.76888f
C315 COMP_2_0.vb.t10 VGND 0.98196f
C316 COMP_2_0.vb.t8 VGND 0.65156f
C317 COMP_2_0.vb.n0 VGND 0.99593f
C318 COMP_2_0.vb.t6 VGND 0.65142f
C319 COMP_2_0.vb.n1 VGND 0.69015f
C320 COMP_2_0.vb.t7 VGND 0.65156f
C321 COMP_2_0.vb.n2 VGND 0.68949f
C322 COMP_2_0.vb.n3 VGND 0.57305f
C323 COMP_2_0.vb.n4 VGND 0.66625f
C324 COMP_2_0.vb.t2 VGND 0.50446f
C325 COMP_2_0.vb.n5 VGND 0.68995f
C326 COMP_2_0.vb.n6 VGND 0.1103f
C327 COMP_2_0.vb.t0 VGND 0.00934f
C328 COMP_2_0.vb.t1 VGND 0.00912f
C329 COMP_2_0.vb.n7 VGND 0.061f
C330 COMP_2_0.vb.n8 VGND 0.05645f
C331 COMP_2_0.vb.t9 VGND 1.61449f
C332 a_11329_22619.n0 VGND 0.01625f
C333 a_11329_22619.t8 VGND 2.45052f
C334 a_11329_22619.n1 VGND 1.00743f
C335 a_11329_22619.t7 VGND 2.48837f
C336 a_11329_22619.n2 VGND 0.0167f
C337 a_11329_22619.t3 VGND 1.24369f
C338 a_11329_22619.t4 VGND 0.01808f
C339 a_11329_22619.n3 VGND 0.04438f
C340 a_11329_22619.n4 VGND 1.08276f
C341 a_11329_22619.n5 VGND 0.05617f
C342 a_11329_22619.n6 VGND 0.97711f
C343 a_11329_22619.n7 VGND 0.07001f
C344 a_11329_22619.t5 VGND 1.22817f
C345 a_11329_22619.n8 VGND 1.15569f
C346 a_11329_22619.t6 VGND 0.01839f
C347 a_11329_22619.n9 VGND 0.09033f
C348 a_11329_22619.t1 VGND 0.14735f
C349 a_11329_22619.t2 VGND 0.07693f
C350 a_11329_22619.n10 VGND 1.1393f
C351 a_11329_22619.n11 VGND 0.21407f
C352 a_11329_22619.n12 VGND 0.55062f
C353 a_11329_22619.t0 VGND 0.00771f
C354 delay_1_0.vd_n.t6 VGND 3.75842f
C355 delay_1_0.vd_n.t4 VGND 1.90817f
C356 delay_1_0.vd_n.n0 VGND 1.33579f
C357 delay_1_0.vd_n.t3 VGND 3.75854f
C358 delay_1_0.vd_n.t2 VGND 1.90817f
C359 delay_1_0.vd_n.n1 VGND 1.8782f
C360 delay_1_0.vd_n.n2 VGND 0.64982f
C361 delay_1_0.vd_n.t0 VGND 0
C362 delay_1_0.vd_n.n3 VGND 0.00897f
C363 delay_1_0.vd_n.t1 VGND 0.04603f
C364 delay_1_0.vd_n.t5 VGND 0.04464f
C365 delay_1_0.vd_n.n4 VGND 0.12629f
C366 a_6061_11160.t3 VGND 0.09573f
C367 a_6061_11160.t4 VGND 0.11049f
C368 a_6061_11160.t0 VGND 0.09572f
C369 a_6061_11160.n0 VGND 1.76398f
C370 a_6061_11160.t2 VGND 0.09572f
C371 a_6061_11160.n1 VGND 0.54262f
C372 a_6061_11160.t1 VGND 0.09573f
C373 COMP_2_0.vin_n.t0 VGND 0.00508f
C374 COMP_2_0.vin_n.t1 VGND 0.00501f
C375 COMP_2_0.vin_n.n0 VGND 0.04201f
C376 COMP_2_0.vin_n.t2 VGND 0.25753f
C377 COMP_2_0.vin_n.t3 VGND 0.24546f
C378 COMP_2_0.vin_n.n1 VGND 0.53438f
C379 a_20802_14722.t1 VGND 4.80071f
C380 a_20802_14722.t3 VGND 4.77949f
C381 a_20802_14722.n0 VGND 0.61852f
C382 a_20802_14722.t2 VGND 0.12764f
C383 a_20802_14722.n1 VGND 0.07316f
C384 a_20802_14722.t0 VGND 0
C385 a_5453_6767.t1 VGND 0.04355f
C386 a_5453_6767.t10 VGND 0.23632f
C387 a_5453_6767.n0 VGND 0.4007f
C388 a_5453_6767.t9 VGND 0.65036f
C389 a_5453_6767.t6 VGND 0.53693f
C390 a_5453_6767.n1 VGND 0.40314f
C391 a_5453_6767.t7 VGND 0.01577f
C392 a_5453_6767.n2 VGND 0.04211f
C393 a_5453_6767.n3 VGND 0.044f
C394 a_5453_6767.n4 VGND 0.43346f
C395 a_5453_6767.t3 VGND 0.0286f
C396 a_5453_6767.t2 VGND 0.0207f
C397 a_5453_6767.n5 VGND 0.53447f
C398 a_5453_6767.n6 VGND 0.21427f
C399 a_5453_6767.n7 VGND 0.40078f
C400 a_5453_6767.t8 VGND 0.65036f
C401 a_5453_6767.t4 VGND 0.53693f
C402 a_5453_6767.n8 VGND 0.40315f
C403 a_5453_6767.t5 VGND 0.01577f
C404 a_5453_6767.n9 VGND 0.04222f
C405 a_5453_6767.n10 VGND 0.04309f
C406 a_5453_6767.n11 VGND 0.25782f
C407 a_5453_6767.n12 VGND 0.79698f
C408 a_5453_6767.t0 VGND 0.04852f
C409 latch_sch_0.R.t4 VGND 0.21283f
C410 latch_sch_0.R.t3 VGND 0.13884f
C411 latch_sch_0.R.t1 VGND 0.06845f
C412 latch_sch_0.R.t2 VGND 0.06041f
C413 latch_sch_0.R.n0 VGND 0.77188f
C414 latch_sch_0.R.t0 VGND 0.02593f
C415 latch_sch_0.R.n1 VGND 0.16962f
C416 a_5453_6051.t6 VGND 0.03201f
C417 a_5453_6051.t7 VGND 0.02834f
C418 a_5453_6051.n0 VGND 0.50031f
C419 a_5453_6051.t5 VGND 0.012f
C420 a_5453_6051.n1 VGND 0.20387f
C421 a_5453_6051.t8 VGND 0.1462f
C422 a_5453_6051.n2 VGND 0.25217f
C423 a_5453_6051.t9 VGND 0.40929f
C424 a_5453_6051.t1 VGND 0.3379f
C425 a_5453_6051.n3 VGND 0.25371f
C426 a_5453_6051.t2 VGND 0.00992f
C427 a_5453_6051.n4 VGND 0.0265f
C428 a_5453_6051.n5 VGND 0.02532f
C429 a_5453_6051.n6 VGND 0.36149f
C430 a_5453_6051.n7 VGND 0.25217f
C431 a_5453_6051.t10 VGND 0.40929f
C432 a_5453_6051.t3 VGND 0.3379f
C433 a_5453_6051.n8 VGND 0.25371f
C434 a_5453_6051.t4 VGND 0.00992f
C435 a_5453_6051.n9 VGND 0.0265f
C436 a_5453_6051.n10 VGND 0.02188f
C437 a_5453_6051.n11 VGND 0.11157f
C438 a_5453_6051.n12 VGND 0.26524f
C439 a_5453_6051.t0 VGND 0.01278f
C440 ua[0].t5 VGND 0.08266f
C441 ua[0].t4 VGND 0.08266f
C442 ua[0].n0 VGND 0.20006f
C443 ua[0].t3 VGND 0.08266f
C444 ua[0].t2 VGND 0.08266f
C445 ua[0].n1 VGND 0.20006f
C446 ua[0].t0 VGND 0.08266f
C447 ua[0].t7 VGND 0.08266f
C448 ua[0].n2 VGND 0.21044f
C449 ua[0].n3 VGND 1.59483f
C450 ua[0].n4 VGND 0.85485f
C451 ua[0].t1 VGND 0.08266f
C452 ua[0].t6 VGND 0.08266f
C453 ua[0].n5 VGND 0.20076f
C454 ua[0].n6 VGND 0.84675f
C455 a_21737_7899.t2 VGND 0.04927f
C456 a_21737_7899.n0 VGND 0.08648f
C457 a_21737_7899.n1 VGND 0.10387f
C458 a_21737_7899.n2 VGND 0.10387f
C459 a_21737_7899.n3 VGND 0.10387f
C460 a_21737_7899.t4 VGND 0.27118f
C461 a_21737_7899.t10 VGND 4.17325f
C462 a_21737_7899.n4 VGND 4.82646f
C463 a_21737_7899.n5 VGND 0.10352f
C464 a_21737_7899.t9 VGND 0.27094f
C465 a_21737_7899.n6 VGND 0.20576f
C466 a_21737_7899.t6 VGND 0.27094f
C467 a_21737_7899.n7 VGND 0.10387f
C468 a_21737_7899.n8 VGND 0.10387f
C469 a_21737_7899.t5 VGND 0.27094f
C470 a_21737_7899.n9 VGND 0.10387f
C471 a_21737_7899.t8 VGND 0.27094f
C472 a_21737_7899.n10 VGND 0.10387f
C473 a_21737_7899.n11 VGND 0.10387f
C474 a_21737_7899.t7 VGND 0.27094f
C475 a_21737_7899.n12 VGND 0.10387f
C476 a_21737_7899.t3 VGND 0.27094f
C477 a_21737_7899.n13 VGND 0.20597f
C478 a_21737_7899.t11 VGND 0.27118f
C479 a_21737_7899.n14 VGND 0.1139f
C480 a_21737_7899.t1 VGND 0.15822f
C481 a_21737_7899.n15 VGND 0.0937f
C482 a_21737_7899.n16 VGND 0.14287f
C483 a_21737_7899.n17 VGND 0.31366f
C484 a_21737_7899.t0 VGND 0.22407f
C485 latch_sch_0.Qn.t0 VGND 0.04597f
C486 latch_sch_0.Qn.t1 VGND 0.00676f
C487 latch_sch_0.Qn.t3 VGND 0.00689f
C488 latch_sch_0.Qn.t2 VGND 0.00736f
C489 latch_sch_0.Qn.n0 VGND 0.05385f
C490 latch_sch_0.Qn.t4 VGND 0.01991f
C491 latch_sch_0.Qn.t5 VGND 0.02056f
C492 latch_sch_0.Qn.n1 VGND 0.05871f
C493 latch_sch_0.Qn.n2 VGND 0.01822f
C494 latch_sch_0.Qn.n3 VGND 0.02947f
C495 a_10404_14647.t2 VGND 0.08651f
C496 a_10404_14647.t4 VGND 0.08447f
C497 a_10404_14647.n0 VGND 0.63297f
C498 a_10404_14647.t8 VGND 0.16876f
C499 a_10404_14647.n1 VGND 0.8149f
C500 a_10404_14647.t9 VGND 0.02892f
C501 a_10404_14647.t1 VGND 0.02871f
C502 a_10404_14647.n2 VGND 1.49302f
C503 a_10404_14647.t5 VGND 0.55248f
C504 a_10404_14647.t7 VGND 0.55248f
C505 a_10404_14647.n3 VGND 4.13746f
C506 a_10404_14647.t3 VGND 0.55248f
C507 a_10404_14647.t6 VGND 0.55248f
C508 a_10404_14647.n4 VGND 4.02251f
C509 a_10404_14647.n5 VGND 2.64013f
C510 a_10404_14647.n6 VGND 1.59538f
C511 a_10404_14647.t0 VGND 0.05634f
C512 a_6404_16954.t1 VGND 0.14794f
C513 a_6404_16954.n0 VGND 0.77905f
C514 a_6404_16954.n1 VGND 3.62123f
C515 a_6404_16954.n2 VGND 3.5173f
C516 a_6404_16954.t7 VGND 5.44967f
C517 a_6404_16954.t9 VGND 1.55601f
C518 a_6404_16954.t8 VGND 1.55601f
C519 a_6404_16954.n3 VGND 4.03755f
C520 a_6404_16954.t10 VGND 2.87614f
C521 a_6404_16954.n4 VGND 5.4777f
C522 a_6404_16954.n5 VGND 3.74605f
C523 a_6404_16954.t6 VGND 5.44967f
C524 a_6404_16954.n6 VGND 4.81675f
C525 a_6404_16954.t5 VGND 0.11473f
C526 a_6404_16954.n7 VGND 0.16453f
C527 a_6404_16954.t4 VGND 5.44967f
C528 a_6404_16954.n8 VGND 3.64676f
C529 a_6404_16954.n9 VGND 1.36067f
C530 a_6404_16954.n10 VGND 1.99681f
C531 a_6404_16954.t2 VGND 5.44967f
C532 a_6404_16954.n11 VGND 4.96673f
C533 a_6404_16954.n12 VGND 1.3508f
C534 a_6404_16954.n13 VGND 1.94937f
C535 a_6404_16954.t3 VGND 0.11473f
C536 a_6404_16954.n14 VGND 0.19695f
C537 a_6404_16954.n15 VGND 0.15023f
C538 a_6404_16954.n16 VGND 1.10222f
C539 a_6404_16954.n17 VGND 0.94546f
C540 a_6404_16954.t0 VGND 0.10963f
C541 VCR_0.VT.t10 VGND 0.22493f
C542 VCR_0.VT.t6 VGND 0.02212f
C543 VCR_0.VT.t5 VGND 0.02212f
C544 VCR_0.VT.n0 VGND 0.06478f
C545 VCR_0.VT.t4 VGND 0.02212f
C546 VCR_0.VT.t3 VGND 0.02212f
C547 VCR_0.VT.n1 VGND 0.06478f
C548 VCR_0.VT.t8 VGND 0.02212f
C549 VCR_0.VT.t0 VGND 0.02212f
C550 VCR_0.VT.n2 VGND 0.06478f
C551 VCR_0.VT.t2 VGND 0.02212f
C552 VCR_0.VT.t1 VGND 0.02212f
C553 VCR_0.VT.n3 VGND 0.07261f
C554 VCR_0.VT.n4 VGND 0.3204f
C555 VCR_0.VT.t7 VGND 0.02212f
C556 VCR_0.VT.t9 VGND 0.02212f
C557 VCR_0.VT.n5 VGND 0.06478f
C558 VCR_0.VT.n6 VGND 0.17685f
C559 VCR_0.VT.n7 VGND 0.17685f
C560 VCR_0.VT.n8 VGND 0.17916f
C561 VCR_0.VT.n9 VGND 0.38391f
C562 VCR_0.VT.t11 VGND 0.43289f
C563 VCR_0.VT.t12 VGND 0.41161f
C564 VCR_0.VT.n10 VGND 0.92643f
C565 ua[2].t0 VGND 0.01646f
C566 ua[2].t1 VGND 0.01965f
C567 ua[2].n0 VGND 0.37342f
C568 ua[2].n1 VGND 0.16791f
C569 ua[2].n2 VGND 0.16749f
C570 ua[2].n3 VGND 0.16785f
C571 ua[2].n4 VGND 0.16795f
C572 ua[2].t5 VGND 0.22216f
C573 ua[2].n5 VGND 0.12567f
C574 ua[2].n6 VGND 0.26581f
C575 ua[2].t6 VGND 0.22181f
C576 ua[2].n7 VGND 0.26581f
C577 ua[2].t7 VGND 0.22181f
C578 ua[2].n9 VGND 0.16795f
C579 ua[2].n10 VGND 0.16775f
C580 ua[2].t8 VGND 0.22181f
C581 ua[2].n12 VGND 0.16775f
C582 ua[2].t4 VGND 0.22181f
C583 ua[2].n14 VGND 0.16785f
C584 ua[2].n15 VGND 0.16766f
C585 ua[2].t2 VGND 0.22181f
C586 ua[2].n17 VGND 0.16766f
C587 ua[2].t3 VGND 0.22181f
C588 ua[2].n19 VGND 0.16749f
C589 ua[2].n20 VGND 0.16775f
C590 ua[2].t11 VGND 0.22181f
C591 ua[2].n22 VGND 0.16775f
C592 ua[2].t9 VGND 0.22181f
C593 ua[2].n24 VGND 0.26379f
C594 ua[2].t10 VGND 0.22181f
C595 ua[2].n25 VGND 0.06516f
C596 ua[2].n26 VGND 0.1733f
C597 ua[2].n27 VGND 0.44853f
C598 ua[2].n28 VGND 0.29775f
C599 Timming_0.Vd.t24 VGND 0.04762f
C600 Timming_0.Vd.t1 VGND 0.05163f
C601 Timming_0.Vd.t25 VGND 0.0487f
C602 Timming_0.Vd.n0 VGND 0.37383f
C603 Timming_0.Vd.t27 VGND 0.1403f
C604 Timming_0.Vd.t26 VGND 0.1466f
C605 Timming_0.Vd.n1 VGND 0.50581f
C606 Timming_0.Vd.n2 VGND 0.18145f
C607 Timming_0.Vd.n3 VGND 0.18785f
C608 Timming_0.Vd.t17 VGND 0.12574f
C609 Timming_0.Vd.t3 VGND 0.12574f
C610 Timming_0.Vd.n4 VGND 0.44978f
C611 Timming_0.Vd.t8 VGND 0.12574f
C612 Timming_0.Vd.t15 VGND 0.12574f
C613 Timming_0.Vd.n5 VGND 0.44978f
C614 Timming_0.Vd.t19 VGND 0.12574f
C615 Timming_0.Vd.t22 VGND 0.12574f
C616 Timming_0.Vd.n6 VGND 0.44978f
C617 Timming_0.Vd.t11 VGND 0.12574f
C618 Timming_0.Vd.t23 VGND 0.12574f
C619 Timming_0.Vd.n7 VGND 0.44978f
C620 Timming_0.Vd.t12 VGND 0.12574f
C621 Timming_0.Vd.t10 VGND 0.12574f
C622 Timming_0.Vd.n8 VGND 0.44978f
C623 Timming_0.Vd.t18 VGND 0.12574f
C624 Timming_0.Vd.t5 VGND 0.12574f
C625 Timming_0.Vd.n9 VGND 0.44978f
C626 Timming_0.Vd.t9 VGND 0.12574f
C627 Timming_0.Vd.t6 VGND 0.12574f
C628 Timming_0.Vd.n10 VGND 0.44979f
C629 Timming_0.Vd.t4 VGND 0.12574f
C630 Timming_0.Vd.t16 VGND 0.12574f
C631 Timming_0.Vd.n11 VGND 0.44978f
C632 Timming_0.Vd.t21 VGND 0.12574f
C633 Timming_0.Vd.t2 VGND 0.12574f
C634 Timming_0.Vd.n12 VGND 0.44978f
C635 Timming_0.Vd.t14 VGND 0.12574f
C636 Timming_0.Vd.t20 VGND 0.12574f
C637 Timming_0.Vd.n13 VGND 0.44978f
C638 Timming_0.Vd.t7 VGND 0.12574f
C639 Timming_0.Vd.t13 VGND 0.12574f
C640 Timming_0.Vd.n14 VGND 0.44978f
C641 Timming_0.Vd.t0 VGND 0.76395f
C642 Timming_0.Vd.n15 VGND 2.39434f
C643 Timming_0.Vd.n16 VGND 0.78729f
C644 Timming_0.Vd.n17 VGND 0.78729f
C645 Timming_0.Vd.n18 VGND 0.78729f
C646 Timming_0.Vd.n19 VGND 0.78723f
C647 Timming_0.Vd.n20 VGND 0.78729f
C648 Timming_0.Vd.n21 VGND 0.78729f
C649 Timming_0.Vd.n22 VGND 0.78729f
C650 Timming_0.Vd.n23 VGND 0.78729f
C651 Timming_0.Vd.n24 VGND 0.78729f
C652 Timming_0.Vd.n25 VGND 0.87339f
C653 a_16597_7688.t43 VGND 0.08239f
C654 a_16597_7688.n0 VGND 0.07776f
C655 a_16597_7688.n1 VGND 0.03056f
C656 a_16597_7688.t41 VGND 0.28878f
C657 a_16597_7688.n2 VGND 0.35653f
C658 a_16597_7688.n3 VGND 0.14591f
C659 a_16597_7688.t42 VGND 0.37671f
C660 a_16597_7688.n4 VGND 0.14591f
C661 a_16597_7688.n5 VGND 0.21614f
C662 a_16597_7688.t40 VGND 0.37671f
C663 a_16597_7688.n6 VGND 0.16537f
C664 a_16597_7688.n7 VGND 0.13649f
C665 a_16597_7688.n8 VGND 0.10225f
C666 a_16597_7688.n9 VGND 0.10225f
C667 a_16597_7688.n10 VGND 0.10225f
C668 a_16597_7688.n11 VGND 0.10225f
C669 a_16597_7688.n12 VGND 0.10225f
C670 a_16597_7688.n13 VGND 0.10225f
C671 a_16597_7688.n14 VGND 0.10225f
C672 a_16597_7688.n15 VGND 0.10225f
C673 a_16597_7688.n16 VGND 0.10225f
C674 a_16597_7688.t9 VGND 0.28878f
C675 a_16597_7688.n17 VGND 0.35653f
C676 a_16597_7688.n18 VGND 0.14591f
C677 a_16597_7688.t37 VGND 0.08239f
C678 a_16597_7688.t11 VGND 0.08239f
C679 a_16597_7688.n19 VGND 0.17473f
C680 a_16597_7688.n20 VGND 0.30041f
C681 a_16597_7688.n21 VGND 0.14591f
C682 a_16597_7688.n22 VGND 0.14591f
C683 a_16597_7688.t19 VGND 0.08239f
C684 a_16597_7688.t39 VGND 0.08239f
C685 a_16597_7688.n23 VGND 0.17473f
C686 a_16597_7688.n24 VGND 0.30041f
C687 a_16597_7688.n25 VGND 0.14591f
C688 a_16597_7688.n26 VGND 0.14591f
C689 a_16597_7688.t27 VGND 0.08239f
C690 a_16597_7688.t31 VGND 0.08239f
C691 a_16597_7688.n27 VGND 0.17473f
C692 a_16597_7688.n28 VGND 0.30041f
C693 a_16597_7688.n29 VGND 0.14591f
C694 a_16597_7688.n30 VGND 0.14591f
C695 a_16597_7688.t15 VGND 0.08239f
C696 a_16597_7688.t17 VGND 0.08239f
C697 a_16597_7688.n31 VGND 0.17473f
C698 a_16597_7688.n32 VGND 0.30041f
C699 a_16597_7688.n33 VGND 0.14591f
C700 a_16597_7688.n34 VGND 0.14591f
C701 a_16597_7688.t7 VGND 0.08239f
C702 a_16597_7688.t35 VGND 0.08239f
C703 a_16597_7688.n35 VGND 0.17473f
C704 a_16597_7688.n36 VGND 0.30041f
C705 a_16597_7688.n37 VGND 0.14591f
C706 a_16597_7688.t0 VGND 0.37671f
C707 a_16597_7688.n38 VGND 0.14591f
C708 a_16597_7688.n39 VGND 0.03056f
C709 a_16597_7688.n40 VGND 0.14591f
C710 a_16597_7688.t6 VGND 0.37671f
C711 a_16597_7688.n41 VGND 0.14591f
C712 a_16597_7688.n42 VGND 0.07776f
C713 a_16597_7688.t34 VGND 0.37671f
C714 a_16597_7688.n43 VGND 0.14591f
C715 a_16597_7688.t21 VGND 0.08239f
C716 a_16597_7688.t13 VGND 0.08239f
C717 a_16597_7688.n44 VGND 0.17473f
C718 a_16597_7688.n45 VGND 0.30041f
C719 a_16597_7688.n46 VGND 0.07776f
C720 a_16597_7688.n47 VGND 0.14591f
C721 a_16597_7688.t20 VGND 0.37671f
C722 a_16597_7688.n48 VGND 0.14591f
C723 a_16597_7688.n49 VGND 0.03056f
C724 a_16597_7688.t12 VGND 0.37671f
C725 a_16597_7688.n50 VGND 0.14591f
C726 a_16597_7688.n51 VGND 0.03056f
C727 a_16597_7688.n52 VGND 0.14591f
C728 a_16597_7688.t14 VGND 0.37671f
C729 a_16597_7688.n53 VGND 0.14591f
C730 a_16597_7688.n54 VGND 0.07776f
C731 a_16597_7688.t16 VGND 0.37671f
C732 a_16597_7688.n55 VGND 0.14591f
C733 a_16597_7688.t23 VGND 0.08239f
C734 a_16597_7688.t3 VGND 0.08239f
C735 a_16597_7688.n56 VGND 0.17473f
C736 a_16597_7688.n57 VGND 0.30041f
C737 a_16597_7688.n58 VGND 0.07776f
C738 a_16597_7688.n59 VGND 0.14591f
C739 a_16597_7688.t22 VGND 0.37671f
C740 a_16597_7688.n60 VGND 0.14591f
C741 a_16597_7688.n61 VGND 0.03056f
C742 a_16597_7688.t2 VGND 0.37671f
C743 a_16597_7688.n62 VGND 0.14591f
C744 a_16597_7688.n63 VGND 0.03056f
C745 a_16597_7688.n64 VGND 0.14591f
C746 a_16597_7688.t26 VGND 0.37671f
C747 a_16597_7688.n65 VGND 0.14591f
C748 a_16597_7688.n66 VGND 0.07776f
C749 a_16597_7688.t30 VGND 0.37671f
C750 a_16597_7688.n67 VGND 0.14591f
C751 a_16597_7688.t33 VGND 0.08239f
C752 a_16597_7688.t29 VGND 0.08239f
C753 a_16597_7688.n68 VGND 0.17473f
C754 a_16597_7688.n69 VGND 0.30041f
C755 a_16597_7688.n70 VGND 0.07776f
C756 a_16597_7688.n71 VGND 0.14591f
C757 a_16597_7688.t32 VGND 0.37671f
C758 a_16597_7688.n72 VGND 0.14591f
C759 a_16597_7688.n73 VGND 0.03056f
C760 a_16597_7688.t28 VGND 0.37671f
C761 a_16597_7688.n74 VGND 0.14591f
C762 a_16597_7688.n75 VGND 0.03056f
C763 a_16597_7688.n76 VGND 0.14591f
C764 a_16597_7688.t18 VGND 0.37671f
C765 a_16597_7688.n77 VGND 0.14591f
C766 a_16597_7688.n78 VGND 0.07776f
C767 a_16597_7688.t38 VGND 0.37671f
C768 a_16597_7688.n79 VGND 0.14591f
C769 a_16597_7688.t25 VGND 0.08239f
C770 a_16597_7688.t5 VGND 0.08239f
C771 a_16597_7688.n80 VGND 0.17473f
C772 a_16597_7688.n81 VGND 0.30041f
C773 a_16597_7688.n82 VGND 0.07776f
C774 a_16597_7688.n83 VGND 0.14591f
C775 a_16597_7688.t24 VGND 0.37671f
C776 a_16597_7688.n84 VGND 0.14591f
C777 a_16597_7688.n85 VGND 0.03056f
C778 a_16597_7688.t4 VGND 0.37671f
C779 a_16597_7688.n86 VGND 0.14591f
C780 a_16597_7688.n87 VGND 0.03056f
C781 a_16597_7688.n88 VGND 0.14591f
C782 a_16597_7688.t36 VGND 0.37671f
C783 a_16597_7688.n89 VGND 0.14591f
C784 a_16597_7688.n90 VGND 0.07776f
C785 a_16597_7688.t10 VGND 0.37671f
C786 a_16597_7688.n91 VGND 0.14591f
C787 a_16597_7688.n92 VGND 0.21614f
C788 a_16597_7688.t8 VGND 0.37671f
C789 a_16597_7688.n93 VGND 0.16537f
C790 a_16597_7688.n94 VGND 0.1112f
C791 a_16597_7688.t44 VGND 0.0328f
C792 a_16597_7688.n95 VGND 0.28522f
C793 a_16597_7688.n96 VGND 0.15707f
C794 a_16597_7688.n97 VGND 0.15707f
C795 a_16597_7688.n98 VGND 0.15707f
C796 a_16597_7688.n99 VGND 0.15707f
C797 a_16597_7688.n100 VGND 0.15707f
C798 a_16597_7688.n101 VGND 0.15707f
C799 a_16597_7688.n102 VGND 0.15707f
C800 a_16597_7688.n103 VGND 0.15707f
C801 a_16597_7688.n104 VGND 0.15707f
C802 a_16597_7688.n105 VGND 0.23784f
C803 a_16597_7688.n106 VGND 0.10225f
C804 a_16597_7688.n107 VGND 0.30041f
C805 a_16597_7688.n108 VGND 0.17473f
C806 a_16597_7688.t1 VGND 0.08239f
C807 VAPWR.n0 VGND 0.26446f
C808 VAPWR.t25 VGND 0.00799f
C809 VAPWR.n1 VGND 0.33238f
C810 VAPWR.n2 VGND 0.1954f
C811 VAPWR.n3 VGND 0.27614f
C812 VAPWR.n4 VGND 0.16119f
C813 VAPWR.n5 VGND 0.0908f
C814 VAPWR.n6 VGND 0.10312f
C815 VAPWR.t28 VGND 0.82964f
C816 VAPWR.n7 VGND 1.50704f
C817 VAPWR.n8 VGND 0.07254f
C818 VAPWR.n9 VGND 0.26056f
C819 VAPWR.n10 VGND 0.03574f
C820 VAPWR.n11 VGND 0.25486f
C821 VAPWR.n12 VGND 0.2099f
C822 VAPWR.n13 VGND 0.23129f
C823 VAPWR.n14 VGND 0.00481f
C824 VAPWR.n15 VGND 0.02008f
C825 VAPWR.n16 VGND 0.04795f
C826 VAPWR.n17 VGND 0.22787f
C827 VAPWR.n18 VGND 0.12504f
C828 VAPWR.n19 VGND 0.10167f
C829 VAPWR.n20 VGND 0.11354f
C830 VAPWR.t0 VGND 0.86676f
C831 VAPWR.n21 VGND 0.03413f
C832 VAPWR.n22 VGND 0.03419f
C833 VAPWR.n23 VGND 0.03419f
C834 VAPWR.n24 VGND 0.0086f
C835 VAPWR.n25 VGND 0.05863f
C836 VAPWR.n26 VGND 0.24024f
C837 VAPWR.n27 VGND 0.06367f
C838 VAPWR.n28 VGND 0.03343f
C839 VAPWR.n29 VGND 0.13802f
C840 VAPWR.n30 VGND 0.03419f
C841 VAPWR.n31 VGND 0.57318f
C842 VAPWR.n32 VGND 0.07104f
C843 VAPWR.n33 VGND 0.10976f
C844 VAPWR.n34 VGND 0.03413f
C845 VAPWR.n35 VGND 0.00842f
C846 VAPWR.n36 VGND 0.0086f
C847 VAPWR.n37 VGND 0.22497f
C848 VAPWR.n38 VGND 0.03413f
C849 VAPWR.n39 VGND 0.03413f
C850 VAPWR.t13 VGND -0.46659f
C851 VAPWR.n40 VGND 0.37237f
C852 VAPWR.n41 VGND 0.63531f
C853 VAPWR.n42 VGND 0.03419f
C854 VAPWR.n43 VGND 0.03419f
C855 VAPWR.n44 VGND 0.03413f
C856 VAPWR.n45 VGND 0.07104f
C857 VAPWR.n46 VGND 0.08598f
C858 VAPWR.n47 VGND 0.2003f
C859 VAPWR.n48 VGND 0.05192f
C860 VAPWR.n49 VGND 0.16574f
C861 VAPWR.n50 VGND 0.1192f
C862 VAPWR.n51 VGND 0.09618f
C863 VAPWR.n52 VGND 0.18201f
C864 VAPWR.n53 VGND 0.09339f
C865 VAPWR.n54 VGND 0.19654f
C866 VAPWR.n55 VGND 0.20825f
C867 VAPWR.n56 VGND 0.01673f
C868 VAPWR.n57 VGND 0.1337f
C869 VAPWR.n58 VGND 0.03419f
C870 VAPWR.n59 VGND 0.03413f
C871 VAPWR.n60 VGND 0.03419f
C872 VAPWR.n61 VGND 0.03419f
C873 VAPWR.n62 VGND 0.19947f
C874 VAPWR.n63 VGND 0.03511f
C875 VAPWR.n64 VGND 0.05558f
C876 VAPWR.n65 VGND 0.09378f
C877 VAPWR.n66 VGND 0.00382f
C878 VAPWR.n67 VGND 0.47144f
C879 VAPWR.n68 VGND 0.21439f
C880 VAPWR.n69 VGND 0.04543f
C881 VAPWR.n70 VGND 0.04924f
C882 VAPWR.n71 VGND 0.04762f
C883 VAPWR.n72 VGND 0.03419f
C884 VAPWR.n73 VGND 0.03413f
C885 VAPWR.n74 VGND 0.03413f
C886 VAPWR.n76 VGND 0.37461f
C887 VAPWR.n77 VGND 0.03413f
C888 VAPWR.n78 VGND 0.03419f
C889 VAPWR.n79 VGND 0.03413f
C890 VAPWR.n80 VGND 0.03413f
C891 VAPWR.n81 VGND 0.71247f
C892 VAPWR.n82 VGND 0.71247f
C893 VAPWR.n83 VGND 0.05203f
C894 VAPWR.n84 VGND 0.10407f
C895 VAPWR.n85 VGND 0.08763f
C896 VAPWR.n86 VGND 0.13571f
C897 VAPWR.n87 VGND 0.09189f
C898 VAPWR.n88 VGND 0.10333f
C899 VAPWR.n89 VGND 0.09096f
C900 VAPWR.n90 VGND 0.14254f
C901 VAPWR.n91 VGND 0.0516f
C902 VAPWR.n92 VGND 0.03419f
C903 VAPWR.t27 VGND 1.00768f
C904 VAPWR.n94 VGND 0.03419f
C905 VAPWR.n95 VGND 0.07804f
C906 VAPWR.n96 VGND 0.09119f
C907 VAPWR.n97 VGND 0.14824f
C908 VAPWR.n98 VGND 0.11401f
C909 VAPWR.n99 VGND 0.09087f
C910 VAPWR.n100 VGND 0.04969f
C911 VAPWR.n101 VGND 0.04181f
C912 VAPWR.n102 VGND 0.00483f
C913 VAPWR.n103 VGND 0.06728f
C914 VAPWR.n104 VGND 0.0357f
C915 VAPWR.n105 VGND 0.27602f
C916 VAPWR.n106 VGND 0.19487f
C917 VAPWR.n107 VGND 0.03413f
C918 VAPWR.n108 VGND 0.38384f
C919 VAPWR.n109 VGND 0.03413f
C920 VAPWR.n110 VGND 0.03419f
C921 VAPWR.n111 VGND 0.07248f
C922 VAPWR.n112 VGND 0.07214f
C923 VAPWR.n113 VGND 0.01087f
C924 VAPWR.n114 VGND 0.10672f
C925 VAPWR.n115 VGND 0.05241f
C926 VAPWR.n116 VGND 0.15453f
C927 VAPWR.n117 VGND 0.26138f
C928 VAPWR.n118 VGND 0.17426f
C929 VAPWR.n119 VGND 0.05781f
C930 VAPWR.n120 VGND 0.0782f
C931 VAPWR.n121 VGND 0.02958f
C932 VAPWR.n122 VGND 0.22497f
C933 VAPWR.n123 VGND 0.09897f
C934 VAPWR.n124 VGND 0.06977f
C935 VAPWR.n125 VGND 0.03419f
C936 VAPWR.t15 VGND 0.86676f
C937 VAPWR.n126 VGND 0.03419f
C938 VAPWR.n127 VGND 0.00842f
C939 VAPWR.n128 VGND 0.04965f
C940 VAPWR.n129 VGND 0.04965f
C941 VAPWR.n130 VGND 0.06158f
C942 VAPWR.n131 VGND 0.03413f
C943 VAPWR.n132 VGND 0.57318f
C944 VAPWR.n133 VGND 0.03413f
C945 VAPWR.n134 VGND 0.03419f
C946 VAPWR.n135 VGND 0.06334f
C947 VAPWR.n136 VGND 0.04366f
C948 VAPWR.n137 VGND 0.03242f
C949 VAPWR.n138 VGND 0.08109f
C950 VAPWR.n139 VGND 0.23632f
C951 VAPWR.n140 VGND 0.01355f
C952 VAPWR.n141 VGND 0.05215f
C953 VAPWR.n142 VGND 0.09895f
C954 VAPWR.n143 VGND 0.03413f
C955 VAPWR.n144 VGND 0.61508f
C956 VAPWR.n145 VGND 0.20262f
C957 VAPWR.n146 VGND 0.0274f
C958 VAPWR.n147 VGND 0.18198f
C959 VAPWR.n148 VGND 0.34291f
C960 VAPWR.n149 VGND 0.75701f
C961 VAPWR.n150 VGND 0.22792f
C962 VAPWR.n151 VGND 0.0907f
C963 VAPWR.n152 VGND 0.17526f
C964 VAPWR.n153 VGND 0.05802f
C965 VAPWR.t24 VGND 0.37028f
C966 VAPWR.n154 VGND 0.05802f
C967 VAPWR.n155 VGND 0.19376f
C968 VAPWR.n156 VGND 0.0183f
C969 VAPWR.n157 VGND 0.15709f
C970 VAPWR.n158 VGND 0.15822f
C971 VAPWR.n159 VGND 0.42429f
C972 VAPWR.n160 VGND 0.38379f
C973 VAPWR.n161 VGND 0.0484f
C974 VAPWR.n162 VGND 0
C975 VAPWR.n163 VGND 0.0898f
C976 VAPWR.n164 VGND 0.03527f
C977 VAPWR.n165 VGND 0
C978 VAPWR.n166 VGND 0
C979 VAPWR.n167 VGND 0.04275f
C980 VAPWR.n168 VGND 0.04493f
C981 VAPWR.n169 VGND 0.04254f
C982 VAPWR.n170 VGND 0.08383f
C983 VAPWR.n171 VGND 0.09307f
C984 VAPWR.t31 VGND 0.09329f
C985 VAPWR.t36 VGND 0.05804f
C986 VAPWR.t2 VGND 0.09463f
C987 VAPWR.t7 VGND 0.05755f
C988 VAPWR.n172 VGND 0.03482f
C989 VAPWR.n173 VGND 0.01643f
C990 VAPWR.n174 VGND 0.03853f
C991 VAPWR.n175 VGND 0.01643f
C992 VAPWR.n176 VGND 0.07774f
C993 VAPWR.n177 VGND 0.04363f
C994 VAPWR.n178 VGND 0.10756f
C995 VAPWR.t37 VGND 0.002f
C996 VAPWR.t8 VGND 0.002f
C997 VAPWR.n179 VGND 0.00428f
C998 VAPWR.n180 VGND 0.0654f
C999 VAPWR.n181 VGND 0.00217f
C1000 VAPWR.n182 VGND 0.03417f
C1001 VAPWR.n183 VGND 0
C1002 VAPWR.n184 VGND 0.03393f
C1003 VAPWR.n185 VGND 0.01115f
C1004 VAPWR.n186 VGND 0.47523f
C1005 VAPWR.n187 VGND 3.64383f
C1006 VAPWR.n188 VGND 1.51226f
C1007 VAPWR.n189 VGND 0.04955f
C1008 VAPWR.n190 VGND 1.12227f
C1009 VAPWR.n191 VGND 0.25056f
C1010 VAPWR.n192 VGND 0.82544f
C1011 VAPWR.n193 VGND 0.62764f
C1012 VAPWR.n194 VGND 0.05083f
C1013 VAPWR.n195 VGND 0.59468f
C1014 VAPWR.n196 VGND 0.09124f
C1015 VAPWR.n197 VGND 0.11027f
C1016 VAPWR.t3 VGND 7.44756f
C1017 VAPWR.n198 VGND 0.11027f
C1018 VAPWR.n199 VGND 0.00238f
C1019 VAPWR.n200 VGND 0.13263f
C1020 VAPWR.n201 VGND 0.04993f
C1021 VAPWR.n202 VGND 0.0527f
C1022 VAPWR.n203 VGND 0.74593f
C1023 VAPWR.n204 VGND 0.784f
C1024 VAPWR.n205 VGND 0.08527f
C1025 VAPWR.n206 VGND 0.0527f
C1026 VAPWR.n207 VGND 0.1987f
C1027 VAPWR.n208 VGND 0.15274f
C1028 VAPWR.n209 VGND 0.10305f
C1029 VAPWR.n210 VGND 0.00612f
C1030 VAPWR.n211 VGND 0.74593f
C1031 VAPWR.n212 VGND 0.05374f
C1032 VAPWR.t11 VGND 0.82121f
C1033 VAPWR.n214 VGND 0.05374f
C1034 VAPWR.n215 VGND 0.10762f
C1035 VAPWR.n216 VGND 0.12641f
C1036 VAPWR.n217 VGND 0.09334f
C1037 VAPWR.n218 VGND 0.05374f
C1038 VAPWR.t14 VGND 0.82121f
C1039 VAPWR.n220 VGND 0.05374f
C1040 VAPWR.n221 VGND 0.01443f
C1041 VAPWR.n222 VGND 0.0375f
C1042 VAPWR.n223 VGND 0.0125f
C1043 VAPWR.n224 VGND 0.15696f
C1044 VAPWR.n225 VGND 0.01508f
C1045 VAPWR.n226 VGND 0.00929f
C1046 VAPWR.n227 VGND 0.00858f
C1047 VAPWR.n228 VGND 0.2844f
C1048 VAPWR.n229 VGND 0.07842f
C1049 VAPWR.n230 VGND 0.04687f
C1050 VAPWR.n231 VGND 0.04687f
C1051 VAPWR.n232 VGND 0.09124f
C1052 VAPWR.n233 VGND 0.05025f
C1053 VAPWR.n234 VGND 7.44756f
C1054 VAPWR.n235 VGND 0.10986f
C1055 VAPWR.n236 VGND 0.11027f
C1056 VAPWR.n237 VGND 4.05088f
C1057 VAPWR.n238 VGND 0.10986f
C1058 VAPWR.n239 VGND 0.09083f
C1059 VAPWR.n240 VGND 1.03757f
C1060 VAPWR.n241 VGND 0.02752f
C1061 VAPWR.n242 VGND 0.49064f
C1062 VAPWR.n243 VGND 0.11995f
C1063 VAPWR.n244 VGND 0.23974f
C1064 VAPWR.n245 VGND 0.68783f
C1065 VAPWR.n246 VGND 0.0619f
C1066 VAPWR.n247 VGND 1.68654f
C1067 VAPWR.n248 VGND 0.58672f
C1068 VAPWR.n249 VGND 0.68066f
C1069 VAPWR.n250 VGND 0.17917f
C1070 VAPWR.n251 VGND 0.19919f
C1071 VAPWR.n252 VGND 0.63063f
C1072 VAPWR.n253 VGND 0.11731f
C1073 VAPWR.n254 VGND 0.10723f
C1074 VAPWR.n255 VGND 0.10723f
C1075 VAPWR.n256 VGND 2.10244f
C1076 VAPWR.n257 VGND 0.11054f
C1077 VAPWR.n258 VGND 2.10244f
C1078 VAPWR.n259 VGND 0.10574f
C1079 VAPWR.n260 VGND 0.11186f
C1080 VAPWR.n261 VGND 0.11215f
C1081 VAPWR.n262 VGND 0.57892f
C1082 VAPWR.n263 VGND 0.02298f
C1083 VAPWR.n264 VGND 0.04802f
C1084 VAPWR.n265 VGND 0.14943f
C1085 VAPWR.n266 VGND 0.02729f
C1086 VAPWR.n267 VGND 0.26822f
C1087 VAPWR.n268 VGND 0.26336f
C1088 VAPWR.n269 VGND 0.15138f
C1089 VAPWR.n270 VGND 0.30498f
C1090 VAPWR.n271 VGND 0.64903f
C1091 VAPWR.n272 VGND 0.37959f
C1092 VAPWR.n273 VGND 0.70522f
C1093 VAPWR.n274 VGND 0.43033f
C1094 VAPWR.n275 VGND 0.19928f
C1095 VAPWR.n276 VGND 0.29927f
C1096 VAPWR.n277 VGND 0.09083f
C1097 VAPWR.n278 VGND 0.06577f
C1098 VAPWR.n279 VGND 0.13384f
C1099 VAPWR.n280 VGND 1.18224f
C1100 VAPWR.n281 VGND 0.48813f
C1101 VAPWR.n282 VGND 0.34271f
C1102 VAPWR.n283 VGND 0.35152f
C1103 VAPWR.n284 VGND 0.01834f
C1104 VAPWR.n285 VGND 0.20262f
C1105 VAPWR.n286 VGND 0.00999f
C1106 VAPWR.n287 VGND 0.02854f
C1107 VAPWR.n288 VGND 0.14462f
C1108 VAPWR.n289 VGND 0.32563f
C1109 VAPWR.n290 VGND 0.11054f
C1110 VAPWR.t6 VGND 3.86534f
C1111 VAPWR.n291 VGND 0.11036f
C1112 VAPWR.n292 VGND 0.29135f
C1113 VAPWR.n293 VGND 0.42639f
C1114 VAPWR.n294 VGND 1.41098f
C1115 VAPWR.n295 VGND 0.98431f
C1116 VAPWR.n296 VGND 0.55454f
C1117 VAPWR.n297 VGND 0.61902f
C1118 VAPWR.n298 VGND 0.05762f
C1119 VAPWR.n299 VGND 0.53332f
C1120 VAPWR.n300 VGND 0.05762f
C1121 VAPWR.n301 VGND 0.43556f
C1122 VAPWR.t4 VGND 0.64722f
C1123 VAPWR.n304 VGND 0.42083f
C1124 VAPWR.n305 VGND 0
C1125 VAPWR.n306 VGND 0.01938f
C1126 VAPWR.n307 VGND 0.02905f
C1127 VAPWR.t5 VGND 0.00747f
C1128 VAPWR.n308 VGND 0.00131f
C1129 VAPWR.n309 VGND 0.00131f
C1130 VAPWR.n310 VGND 0.0015f
C1131 VAPWR.n311 VGND 1.11336f
C1132 VAPWR.n312 VGND 1.15766f
C1133 VAPWR.n313 VGND 0.06346f
C1134 VAPWR.n314 VGND 0.40651f
C1135 VAPWR.n315 VGND 1.30401f
C1136 VAPWR.n316 VGND 0.21491f
C1137 VAPWR.n317 VGND 0.06142f
C1138 VAPWR.n318 VGND 0.11939f
C1139 VAPWR.n319 VGND 0.45958f
C1140 VAPWR.n320 VGND 0.59099f
C1141 VAPWR.n321 VGND 0.11027f
C1142 VAPWR.t1 VGND 7.44756f
C1143 VAPWR.n322 VGND 0.08643f
C1144 VAPWR.n323 VGND 0.1333f
C1145 VAPWR.n324 VGND 0.08643f
C1146 VAPWR.n325 VGND 0.05032f
C1147 VAPWR.n326 VGND 0.38435f
C1148 VAPWR.n327 VGND 0.55891f
C1149 VAPWR.n328 VGND 0.09083f
C1150 VAPWR.n329 VGND 4.05088f
C1151 VAPWR.n330 VGND 0.09083f
C1152 VAPWR.n331 VGND 0.6403f
C1153 VAPWR.n332 VGND 0.29068f
C1154 VAPWR.n333 VGND 1.19759f
C1155 VAPWR.n334 VGND 1.7251f
C1156 VAPWR.n335 VGND 0.31333f
C1157 VAPWR.n336 VGND 1.14567f
C1158 VAPWR.n337 VGND 0.10946f
C1159 VAPWR.n338 VGND 0.04738f
C1160 VAPWR.n339 VGND 0.09184f
C1161 VAPWR.n340 VGND 0.05779f
C1162 VAPWR.n341 VGND 0.66609f
C1163 VAPWR.n342 VGND 0.34037f
C1164 VAPWR.n343 VGND 0.08121f
C1165 VAPWR.n344 VGND 0.33256f
C1166 VAPWR.n345 VGND 0.19305f
C1167 VAPWR.n346 VGND 0.08905f
C1168 VAPWR.n347 VGND 0.05192f
C1169 VAPWR.n348 VGND 0.05192f
C1170 VAPWR.n349 VGND 0.05214f
C1171 VAPWR.n350 VGND 0.42242f
C1172 VAPWR.n351 VGND 0.18954f
C1173 VAPWR.n352 VGND 0.00102f
C1174 VAPWR.n353 VGND 0.08398f
C1175 VAPWR.n354 VGND 0.19993f
C1176 VAPWR.n355 VGND 0.10354f
C1177 VAPWR.n356 VGND 0.10002f
C1178 VAPWR.n357 VGND 0.19258f
C1179 VAPWR.n358 VGND 0.05214f
C1180 VAPWR.t26 VGND 0.64305f
C1181 VAPWR.n361 VGND 0.05214f
C1182 VAPWR.n362 VGND 0.20031f
C1183 VAPWR.n363 VGND 0.09198f
C1184 VAPWR.n364 VGND 0.09451f
C1185 VAPWR.n365 VGND 0.42241f
C1186 VAPWR.n366 VGND 0.05214f
C1187 VAPWR.t12 VGND 0.64305f
C1188 VAPWR.n367 VGND 0.63615f
C1189 VAPWR.n368 VGND 0.01091f
C1190 VAPWR.n369 VGND 0.00645f
C1191 VAPWR.n370 VGND 0.08632f
C1192 VAPWR.n371 VGND 0.00106f
C1193 VAPWR.n372 VGND 0.18959f
C1194 VAPWR.n373 VGND 0.72348f
C1195 VAPWR.n374 VGND 0.11229f
C1196 VAPWR.n375 VGND 0.29504f
C1197 VAPWR.n376 VGND 11.6778f
C1198 VAPWR.n377 VGND 1.16758f
C1199 VAPWR.n378 VGND 31.1923f
C1200 VAPWR.n379 VGND 2.01025f
C1201 VAPWR.n380 VGND 0.12203f
C1202 VAPWR.n381 VGND 0.00661f
C1203 VAPWR.n382 VGND 0.14034f
C1204 VAPWR.n383 VGND 0.32087f
C1205 VAPWR.n384 VGND 0.09837f
C1206 VAPWR.n385 VGND 0.01722f
C1207 VAPWR.n386 VGND 0.12861f
C1208 VAPWR.n387 VGND 0.10127f
C1209 VAPWR.t30 VGND 0.03008f
C1210 VAPWR.t19 VGND 0.06717f
C1211 VAPWR.n388 VGND 0.12945f
C1212 VAPWR.t17 VGND 0.06871f
C1213 VAPWR.t21 VGND 0.01698f
C1214 VAPWR.t35 VGND 0.01698f
C1215 VAPWR.n389 VGND 0.04129f
C1216 VAPWR.t33 VGND 0.01698f
C1217 VAPWR.t23 VGND 0.01698f
C1218 VAPWR.n390 VGND 0.04129f
C1219 VAPWR.t10 VGND 0.01698f
C1220 VAPWR.t39 VGND 0.01698f
C1221 VAPWR.n391 VGND 0.04129f
C1222 VAPWR.n392 VGND 0.18619f
C1223 VAPWR.n393 VGND 0.17016f
C1224 VAPWR.n394 VGND 0.17016f
C1225 VAPWR.n395 VGND 0.1568f
C1226 VAPWR.n396 VGND 0.47735f
C1227 VAPWR.n397 VGND 0.14555f
C1228 VAPWR.n398 VGND 0.52702f
C1229 VAPWR.n399 VGND 0.1587f
C1230 VAPWR.n400 VGND 0.08867f
C1231 VAPWR.n401 VGND 0.42681f
C1232 VAPWR.n403 VGND 0.21926f
C1233 VAPWR.n404 VGND 0.03405f
C1234 VAPWR.n405 VGND 0.03405f
C1235 VAPWR.n406 VGND 0.09221f
C1236 VAPWR.n407 VGND 0.01838f
C1237 VAPWR.n408 VGND 0.02743f
C1238 VAPWR.n409 VGND 0.20199f
C1239 VAPWR.n410 VGND 0.02273f
C1240 VAPWR.n411 VGND 0.03529f
C1241 VAPWR.n412 VGND 0.03267f
C1242 VAPWR.n413 VGND 0.14313f
C1243 VAPWR.n414 VGND 0.03018f
C1244 VAPWR.n415 VGND 0.02228f
C1245 VAPWR.n416 VGND 0.00188f
C1246 VAPWR.n417 VGND 0.01124f
C1247 VAPWR.n418 VGND 0.02992f
C1248 VAPWR.n419 VGND 0.03453f
C1249 VAPWR.n420 VGND 0.03875f
C1250 VAPWR.n421 VGND 0.06123f
C1251 VAPWR.n422 VGND 0.22021f
C1252 VAPWR.n423 VGND 0.06275f
C1253 VAPWR.n424 VGND 0.21926f
C1254 VAPWR.t29 VGND 0.38469f
C1255 VAPWR.n426 VGND 0.28288f
C1256 VAPWR.t18 VGND 0.41168f
C1257 VAPWR.t9 VGND 0.40773f
C1258 VAPWR.t38 VGND 0.40773f
C1259 VAPWR.t32 VGND 0.3058f
C1260 VAPWR.t16 VGND 0.43149f
C1261 VAPWR.t34 VGND 0.40773f
C1262 VAPWR.t20 VGND 0.40773f
C1263 VAPWR.t22 VGND 0.3058f
C1264 VAPWR.n427 VGND 0.1596f
C1265 VAPWR.n428 VGND 0.08858f
C1266 VAPWR.n429 VGND 0.20387f
C1267 VAPWR.n430 VGND 0.08858f
C1268 VAPWR.n431 VGND 0.33495f
C1269 VAPWR.n432 VGND 0.55025f
C1270 VAPWR.n433 VGND 0.18259f
C1271 VAPWR.n434 VGND 0.14104f
C1272 VAPWR.n435 VGND 0.78961f
C1273 VAPWR.n436 VGND 0.80962f
C1274 VAPWR.n437 VGND 0.2448f
C1275 VAPWR.n438 VGND 0.35382f
C1276 VAPWR.n439 VGND 0.16477f
C1277 VAPWR.n440 VGND 0.03075f
C1278 VAPWR.n441 VGND 0.10528f
C1279 VAPWR.n442 VGND 0.02754f
C1280 VAPWR.n443 VGND 0.03859f
C1281 VAPWR.n444 VGND 0.14905f
C1282 VAPWR.n445 VGND 0.51213f
C1283 VAPWR.n446 VGND 0.12475f
C1284 VAPWR.n447 VGND 0.21495f
C1285 VAPWR.n448 VGND 0.09415f
C1286 VAPWR.n449 VGND 0.11511f
C1287 VAPWR.n450 VGND 0.52452f
C1288 VAPWR.n451 VGND 6.45466f
C1289 a_9577_9007.t1 VGND 0.05445f
C1290 a_9577_9007.t4 VGND 0.14275f
C1291 a_9577_9007.t2 VGND 0.13276f
C1292 a_9577_9007.n0 VGND 0.78577f
C1293 a_9577_9007.t5 VGND 0.14275f
C1294 a_9577_9007.t3 VGND 0.13276f
C1295 a_9577_9007.n1 VGND 0.78577f
C1296 a_9577_9007.n2 VGND 0.26691f
C1297 a_9577_9007.n3 VGND 0.65207f
C1298 a_9577_9007.t0 VGND 0.10399f
C1299 a_9039_8199.n0 VGND 0.32899f
C1300 a_9039_8199.t5 VGND 0.7543f
C1301 a_9039_8199.n1 VGND 0.94403f
C1302 a_9039_8199.t6 VGND 0.74151f
C1303 a_9039_8199.t4 VGND 0.03886f
C1304 a_9039_8199.n2 VGND 0.95123f
C1305 a_9039_8199.n3 VGND 0.08202f
C1306 a_9039_8199.t3 VGND 0.08617f
C1307 a_9039_8199.n4 VGND 0.16895f
C1308 a_9039_8199.t2 VGND 0.73852f
C1309 a_9039_8199.n5 VGND 0.40268f
C1310 a_9039_8199.n6 VGND 0.46973f
C1311 a_9039_8199.n7 VGND 0.12955f
C1312 a_9039_8199.n8 VGND 1.06374f
C1313 a_9039_8199.n9 VGND 0.12252f
C1314 a_9039_8199.t0 VGND 0.73852f
C1315 a_9039_8199.n10 VGND 0.36175f
C1316 a_9039_8199.n11 VGND 0.48112f
C1317 a_9039_8199.n12 VGND 0.10964f
C1318 a_9039_8199.t1 VGND 0.08617f
.ends

