magic
tech sky130A
magscale 1 2
timestamp 1755054771
<< nwell >>
rect 6021 30421 10863 31215
rect 6146 16754 10662 19348
rect 8156 14350 10662 15144
rect 11234 14350 20076 19348
rect 20602 14464 21800 18980
rect 7861 11857 10387 12620
rect 5861 11826 10387 11857
rect 5861 10889 10377 11826
rect 11847 11085 12883 11115
rect 5861 10863 10767 10889
rect 5973 8735 7905 10863
rect 8839 8710 10767 10863
rect 11836 10422 12915 11085
rect 11847 10407 12883 10422
rect 24534 7451 25928 8157
rect 24534 4929 26828 7451
<< pwell >>
rect 2620 30182 5686 42404
rect 7420 27094 13442 28279
rect 7370 26983 13442 27094
rect 7420 24621 13442 26983
rect 13621 28135 14961 28288
rect 13621 27101 13774 28135
rect 14808 27101 14961 28135
rect 13621 26948 14961 27101
rect 14965 28135 16305 28288
rect 14965 27101 15118 28135
rect 16152 27101 16305 28135
rect 14965 26948 16305 27101
rect 16309 28135 17649 28288
rect 16309 27101 16462 28135
rect 17496 27101 17649 28135
rect 16309 26948 17649 27101
rect 13621 26791 14961 26944
rect 13621 25757 13774 26791
rect 14808 25757 14961 26791
rect 13621 25604 14961 25757
rect 14965 26791 16305 26944
rect 14965 25757 15118 26791
rect 16152 25757 16305 26791
rect 14965 25604 16305 25757
rect 16309 26791 17649 26944
rect 16309 25757 16462 26791
rect 17496 25757 17649 26791
rect 16309 25604 17649 25757
rect 13621 25447 14961 25600
rect 13621 24413 13774 25447
rect 14808 24413 14961 25447
rect 10813 24284 10907 24347
rect 5894 19828 10907 24284
rect 13621 24260 14961 24413
rect 14965 25447 16305 25600
rect 14965 24413 15118 25447
rect 16152 24413 16305 25447
rect 14965 24260 16305 24413
rect 16309 25447 17649 25600
rect 16309 24413 16462 25447
rect 17496 24413 17649 25447
rect 16309 24260 17649 24413
rect 15615 23477 20071 23877
rect 11159 22361 20071 23477
rect 11166 21089 20071 22205
rect 11166 20689 15622 21089
rect 10813 19719 10907 19828
rect 11235 9192 13459 9908
rect 5283 5793 8595 8657
rect 8869 7941 9765 8657
rect 9841 7942 10737 8658
rect 13931 2441 16405 10863
rect 16427 7430 20301 9946
rect 16423 4903 18311 7359
rect 16423 2441 18311 4897
rect 18548 2441 19838 6405
rect 21479 3621 23995 8127
rect 21264 1669 24242 3185
rect 24408 1763 26924 4019
<< nbase >>
rect 13774 27101 14808 28135
rect 15118 27101 16152 28135
rect 16462 27101 17496 28135
rect 13774 25757 14808 26791
rect 15118 25757 16152 26791
rect 16462 25757 17496 26791
rect 13774 24413 14808 25447
rect 15118 24413 16152 25447
rect 16462 24413 17496 25447
<< mvnmos >>
rect 6152 20056 6252 24056
rect 6638 20056 6738 24056
rect 7124 20056 7224 24056
rect 7610 20056 7710 24056
rect 8096 20056 8196 24056
rect 8582 20056 8682 24056
rect 9068 20056 9168 24056
rect 9554 20056 9654 24056
rect 10040 20056 10140 24056
rect 10526 20056 10626 24056
rect 11387 22619 15387 23219
rect 15843 22619 19843 23619
rect 11394 20947 15394 21947
rect 15843 21347 19843 21947
rect 11463 9450 11563 9650
rect 12019 9450 12119 9650
rect 12575 9450 12675 9650
rect 13131 9450 13231 9650
rect 5511 8199 6711 8399
rect 7167 8199 8367 8399
rect 9097 8199 9537 8399
rect 10069 8200 10509 8400
rect 5511 7483 6711 7683
rect 7167 7483 8367 7683
rect 5511 6767 6711 6967
rect 7167 6767 8367 6967
rect 16655 7688 16755 9688
rect 16813 7688 16913 9688
rect 16971 7688 17071 9688
rect 17129 7688 17229 9688
rect 17287 7688 17387 9688
rect 17445 7688 17545 9688
rect 17603 7688 17703 9688
rect 17761 7688 17861 9688
rect 17919 7688 18019 9688
rect 18077 7688 18177 9688
rect 18235 7688 18335 9688
rect 18393 7688 18493 9688
rect 18551 7688 18651 9688
rect 18709 7688 18809 9688
rect 18867 7688 18967 9688
rect 19025 7688 19125 9688
rect 19183 7688 19283 9688
rect 19341 7688 19441 9688
rect 19499 7688 19599 9688
rect 19657 7688 19757 9688
rect 19815 7688 19915 9688
rect 19973 7688 20073 9688
rect 5511 6051 6711 6251
rect 7167 6051 8367 6251
rect 21492 1927 21692 2927
rect 21750 1927 21950 2927
rect 22008 1927 22208 2927
rect 22266 1927 22466 2927
rect 22524 1927 22724 2927
rect 22782 1927 22982 2927
rect 23040 1927 23240 2927
rect 23298 1927 23498 2927
rect 23556 1927 23756 2927
rect 23814 1927 24014 2927
<< mvpmos >>
rect 6279 30718 8279 30918
rect 8605 30718 10605 30918
rect 6404 18751 10404 19051
rect 6404 18215 10404 18515
rect 6404 17051 10404 17651
rect 11492 17051 15492 19051
rect 15818 17051 19818 19051
rect 8414 14647 10404 14847
rect 11492 14647 15492 16647
rect 15818 14647 19818 16647
rect 20899 14722 20999 18722
rect 21403 14722 21503 18722
rect 8119 12123 10129 12323
rect 6119 11160 10119 11560
rect 6231 10074 6711 10574
rect 7167 10074 7647 10574
rect 9097 10092 9577 10592
rect 10029 10092 10509 10592
rect 12079 10665 12179 10865
rect 12237 10665 12337 10865
rect 12395 10665 12495 10865
rect 12553 10665 12653 10865
rect 6231 9032 6711 9532
rect 7167 9032 7647 9532
rect 9097 9007 9577 9507
rect 10029 9007 10509 9507
rect 24831 7699 25631 7899
rect 24831 6993 26531 7193
rect 24831 6735 26531 6935
rect 24831 6477 26531 6677
rect 24831 6219 26531 6419
rect 24831 5961 26531 6161
rect 24831 5703 26531 5903
rect 24831 5445 26531 5645
rect 24831 5187 26531 5387
<< mvnnmos >>
rect 16681 5131 16881 7131
rect 17267 5131 17467 7131
rect 17853 5131 18053 7131
rect 16681 2669 16881 4669
rect 17267 2669 17467 4669
rect 17853 2669 18053 4669
rect 21737 6099 23737 7899
rect 21737 3849 23737 5649
rect 24666 1991 26666 3791
<< pdiff >>
rect 13951 27904 14631 27958
rect 13951 27870 14003 27904
rect 14037 27870 14093 27904
rect 14127 27870 14183 27904
rect 14217 27870 14273 27904
rect 14307 27870 14363 27904
rect 14397 27870 14453 27904
rect 14487 27870 14543 27904
rect 14577 27870 14631 27904
rect 13951 27814 14631 27870
rect 13951 27780 14003 27814
rect 14037 27780 14093 27814
rect 14127 27780 14183 27814
rect 14217 27780 14273 27814
rect 14307 27780 14363 27814
rect 14397 27780 14453 27814
rect 14487 27780 14543 27814
rect 14577 27780 14631 27814
rect 13951 27724 14631 27780
rect 13951 27690 14003 27724
rect 14037 27690 14093 27724
rect 14127 27690 14183 27724
rect 14217 27690 14273 27724
rect 14307 27690 14363 27724
rect 14397 27690 14453 27724
rect 14487 27690 14543 27724
rect 14577 27690 14631 27724
rect 13951 27634 14631 27690
rect 13951 27600 14003 27634
rect 14037 27600 14093 27634
rect 14127 27600 14183 27634
rect 14217 27600 14273 27634
rect 14307 27600 14363 27634
rect 14397 27600 14453 27634
rect 14487 27600 14543 27634
rect 14577 27600 14631 27634
rect 13951 27544 14631 27600
rect 13951 27510 14003 27544
rect 14037 27510 14093 27544
rect 14127 27510 14183 27544
rect 14217 27510 14273 27544
rect 14307 27510 14363 27544
rect 14397 27510 14453 27544
rect 14487 27510 14543 27544
rect 14577 27510 14631 27544
rect 13951 27454 14631 27510
rect 13951 27420 14003 27454
rect 14037 27420 14093 27454
rect 14127 27420 14183 27454
rect 14217 27420 14273 27454
rect 14307 27420 14363 27454
rect 14397 27420 14453 27454
rect 14487 27420 14543 27454
rect 14577 27420 14631 27454
rect 13951 27364 14631 27420
rect 13951 27330 14003 27364
rect 14037 27330 14093 27364
rect 14127 27330 14183 27364
rect 14217 27330 14273 27364
rect 14307 27330 14363 27364
rect 14397 27330 14453 27364
rect 14487 27330 14543 27364
rect 14577 27330 14631 27364
rect 13951 27278 14631 27330
rect 15295 27904 15975 27958
rect 15295 27870 15347 27904
rect 15381 27870 15437 27904
rect 15471 27870 15527 27904
rect 15561 27870 15617 27904
rect 15651 27870 15707 27904
rect 15741 27870 15797 27904
rect 15831 27870 15887 27904
rect 15921 27870 15975 27904
rect 15295 27814 15975 27870
rect 15295 27780 15347 27814
rect 15381 27780 15437 27814
rect 15471 27780 15527 27814
rect 15561 27780 15617 27814
rect 15651 27780 15707 27814
rect 15741 27780 15797 27814
rect 15831 27780 15887 27814
rect 15921 27780 15975 27814
rect 15295 27724 15975 27780
rect 15295 27690 15347 27724
rect 15381 27690 15437 27724
rect 15471 27690 15527 27724
rect 15561 27690 15617 27724
rect 15651 27690 15707 27724
rect 15741 27690 15797 27724
rect 15831 27690 15887 27724
rect 15921 27690 15975 27724
rect 15295 27634 15975 27690
rect 15295 27600 15347 27634
rect 15381 27600 15437 27634
rect 15471 27600 15527 27634
rect 15561 27600 15617 27634
rect 15651 27600 15707 27634
rect 15741 27600 15797 27634
rect 15831 27600 15887 27634
rect 15921 27600 15975 27634
rect 15295 27544 15975 27600
rect 15295 27510 15347 27544
rect 15381 27510 15437 27544
rect 15471 27510 15527 27544
rect 15561 27510 15617 27544
rect 15651 27510 15707 27544
rect 15741 27510 15797 27544
rect 15831 27510 15887 27544
rect 15921 27510 15975 27544
rect 15295 27454 15975 27510
rect 15295 27420 15347 27454
rect 15381 27420 15437 27454
rect 15471 27420 15527 27454
rect 15561 27420 15617 27454
rect 15651 27420 15707 27454
rect 15741 27420 15797 27454
rect 15831 27420 15887 27454
rect 15921 27420 15975 27454
rect 15295 27364 15975 27420
rect 15295 27330 15347 27364
rect 15381 27330 15437 27364
rect 15471 27330 15527 27364
rect 15561 27330 15617 27364
rect 15651 27330 15707 27364
rect 15741 27330 15797 27364
rect 15831 27330 15887 27364
rect 15921 27330 15975 27364
rect 15295 27278 15975 27330
rect 16639 27904 17319 27958
rect 16639 27870 16691 27904
rect 16725 27870 16781 27904
rect 16815 27870 16871 27904
rect 16905 27870 16961 27904
rect 16995 27870 17051 27904
rect 17085 27870 17141 27904
rect 17175 27870 17231 27904
rect 17265 27870 17319 27904
rect 16639 27814 17319 27870
rect 16639 27780 16691 27814
rect 16725 27780 16781 27814
rect 16815 27780 16871 27814
rect 16905 27780 16961 27814
rect 16995 27780 17051 27814
rect 17085 27780 17141 27814
rect 17175 27780 17231 27814
rect 17265 27780 17319 27814
rect 16639 27724 17319 27780
rect 16639 27690 16691 27724
rect 16725 27690 16781 27724
rect 16815 27690 16871 27724
rect 16905 27690 16961 27724
rect 16995 27690 17051 27724
rect 17085 27690 17141 27724
rect 17175 27690 17231 27724
rect 17265 27690 17319 27724
rect 16639 27634 17319 27690
rect 16639 27600 16691 27634
rect 16725 27600 16781 27634
rect 16815 27600 16871 27634
rect 16905 27600 16961 27634
rect 16995 27600 17051 27634
rect 17085 27600 17141 27634
rect 17175 27600 17231 27634
rect 17265 27600 17319 27634
rect 16639 27544 17319 27600
rect 16639 27510 16691 27544
rect 16725 27510 16781 27544
rect 16815 27510 16871 27544
rect 16905 27510 16961 27544
rect 16995 27510 17051 27544
rect 17085 27510 17141 27544
rect 17175 27510 17231 27544
rect 17265 27510 17319 27544
rect 16639 27454 17319 27510
rect 16639 27420 16691 27454
rect 16725 27420 16781 27454
rect 16815 27420 16871 27454
rect 16905 27420 16961 27454
rect 16995 27420 17051 27454
rect 17085 27420 17141 27454
rect 17175 27420 17231 27454
rect 17265 27420 17319 27454
rect 16639 27364 17319 27420
rect 16639 27330 16691 27364
rect 16725 27330 16781 27364
rect 16815 27330 16871 27364
rect 16905 27330 16961 27364
rect 16995 27330 17051 27364
rect 17085 27330 17141 27364
rect 17175 27330 17231 27364
rect 17265 27330 17319 27364
rect 16639 27278 17319 27330
rect 13951 26560 14631 26614
rect 13951 26526 14003 26560
rect 14037 26526 14093 26560
rect 14127 26526 14183 26560
rect 14217 26526 14273 26560
rect 14307 26526 14363 26560
rect 14397 26526 14453 26560
rect 14487 26526 14543 26560
rect 14577 26526 14631 26560
rect 13951 26470 14631 26526
rect 13951 26436 14003 26470
rect 14037 26436 14093 26470
rect 14127 26436 14183 26470
rect 14217 26436 14273 26470
rect 14307 26436 14363 26470
rect 14397 26436 14453 26470
rect 14487 26436 14543 26470
rect 14577 26436 14631 26470
rect 13951 26380 14631 26436
rect 13951 26346 14003 26380
rect 14037 26346 14093 26380
rect 14127 26346 14183 26380
rect 14217 26346 14273 26380
rect 14307 26346 14363 26380
rect 14397 26346 14453 26380
rect 14487 26346 14543 26380
rect 14577 26346 14631 26380
rect 13951 26290 14631 26346
rect 13951 26256 14003 26290
rect 14037 26256 14093 26290
rect 14127 26256 14183 26290
rect 14217 26256 14273 26290
rect 14307 26256 14363 26290
rect 14397 26256 14453 26290
rect 14487 26256 14543 26290
rect 14577 26256 14631 26290
rect 13951 26200 14631 26256
rect 13951 26166 14003 26200
rect 14037 26166 14093 26200
rect 14127 26166 14183 26200
rect 14217 26166 14273 26200
rect 14307 26166 14363 26200
rect 14397 26166 14453 26200
rect 14487 26166 14543 26200
rect 14577 26166 14631 26200
rect 13951 26110 14631 26166
rect 13951 26076 14003 26110
rect 14037 26076 14093 26110
rect 14127 26076 14183 26110
rect 14217 26076 14273 26110
rect 14307 26076 14363 26110
rect 14397 26076 14453 26110
rect 14487 26076 14543 26110
rect 14577 26076 14631 26110
rect 13951 26020 14631 26076
rect 13951 25986 14003 26020
rect 14037 25986 14093 26020
rect 14127 25986 14183 26020
rect 14217 25986 14273 26020
rect 14307 25986 14363 26020
rect 14397 25986 14453 26020
rect 14487 25986 14543 26020
rect 14577 25986 14631 26020
rect 13951 25934 14631 25986
rect 15295 26560 15975 26614
rect 15295 26526 15347 26560
rect 15381 26526 15437 26560
rect 15471 26526 15527 26560
rect 15561 26526 15617 26560
rect 15651 26526 15707 26560
rect 15741 26526 15797 26560
rect 15831 26526 15887 26560
rect 15921 26526 15975 26560
rect 15295 26470 15975 26526
rect 15295 26436 15347 26470
rect 15381 26436 15437 26470
rect 15471 26436 15527 26470
rect 15561 26436 15617 26470
rect 15651 26436 15707 26470
rect 15741 26436 15797 26470
rect 15831 26436 15887 26470
rect 15921 26436 15975 26470
rect 15295 26380 15975 26436
rect 15295 26346 15347 26380
rect 15381 26346 15437 26380
rect 15471 26346 15527 26380
rect 15561 26346 15617 26380
rect 15651 26346 15707 26380
rect 15741 26346 15797 26380
rect 15831 26346 15887 26380
rect 15921 26346 15975 26380
rect 15295 26290 15975 26346
rect 15295 26256 15347 26290
rect 15381 26256 15437 26290
rect 15471 26256 15527 26290
rect 15561 26256 15617 26290
rect 15651 26256 15707 26290
rect 15741 26256 15797 26290
rect 15831 26256 15887 26290
rect 15921 26256 15975 26290
rect 15295 26200 15975 26256
rect 15295 26166 15347 26200
rect 15381 26166 15437 26200
rect 15471 26166 15527 26200
rect 15561 26166 15617 26200
rect 15651 26166 15707 26200
rect 15741 26166 15797 26200
rect 15831 26166 15887 26200
rect 15921 26166 15975 26200
rect 15295 26110 15975 26166
rect 15295 26076 15347 26110
rect 15381 26076 15437 26110
rect 15471 26076 15527 26110
rect 15561 26076 15617 26110
rect 15651 26076 15707 26110
rect 15741 26076 15797 26110
rect 15831 26076 15887 26110
rect 15921 26076 15975 26110
rect 15295 26020 15975 26076
rect 15295 25986 15347 26020
rect 15381 25986 15437 26020
rect 15471 25986 15527 26020
rect 15561 25986 15617 26020
rect 15651 25986 15707 26020
rect 15741 25986 15797 26020
rect 15831 25986 15887 26020
rect 15921 25986 15975 26020
rect 15295 25934 15975 25986
rect 16639 26560 17319 26614
rect 16639 26526 16691 26560
rect 16725 26526 16781 26560
rect 16815 26526 16871 26560
rect 16905 26526 16961 26560
rect 16995 26526 17051 26560
rect 17085 26526 17141 26560
rect 17175 26526 17231 26560
rect 17265 26526 17319 26560
rect 16639 26470 17319 26526
rect 16639 26436 16691 26470
rect 16725 26436 16781 26470
rect 16815 26436 16871 26470
rect 16905 26436 16961 26470
rect 16995 26436 17051 26470
rect 17085 26436 17141 26470
rect 17175 26436 17231 26470
rect 17265 26436 17319 26470
rect 16639 26380 17319 26436
rect 16639 26346 16691 26380
rect 16725 26346 16781 26380
rect 16815 26346 16871 26380
rect 16905 26346 16961 26380
rect 16995 26346 17051 26380
rect 17085 26346 17141 26380
rect 17175 26346 17231 26380
rect 17265 26346 17319 26380
rect 16639 26290 17319 26346
rect 16639 26256 16691 26290
rect 16725 26256 16781 26290
rect 16815 26256 16871 26290
rect 16905 26256 16961 26290
rect 16995 26256 17051 26290
rect 17085 26256 17141 26290
rect 17175 26256 17231 26290
rect 17265 26256 17319 26290
rect 16639 26200 17319 26256
rect 16639 26166 16691 26200
rect 16725 26166 16781 26200
rect 16815 26166 16871 26200
rect 16905 26166 16961 26200
rect 16995 26166 17051 26200
rect 17085 26166 17141 26200
rect 17175 26166 17231 26200
rect 17265 26166 17319 26200
rect 16639 26110 17319 26166
rect 16639 26076 16691 26110
rect 16725 26076 16781 26110
rect 16815 26076 16871 26110
rect 16905 26076 16961 26110
rect 16995 26076 17051 26110
rect 17085 26076 17141 26110
rect 17175 26076 17231 26110
rect 17265 26076 17319 26110
rect 16639 26020 17319 26076
rect 16639 25986 16691 26020
rect 16725 25986 16781 26020
rect 16815 25986 16871 26020
rect 16905 25986 16961 26020
rect 16995 25986 17051 26020
rect 17085 25986 17141 26020
rect 17175 25986 17231 26020
rect 17265 25986 17319 26020
rect 16639 25934 17319 25986
rect 13951 25216 14631 25270
rect 13951 25182 14003 25216
rect 14037 25182 14093 25216
rect 14127 25182 14183 25216
rect 14217 25182 14273 25216
rect 14307 25182 14363 25216
rect 14397 25182 14453 25216
rect 14487 25182 14543 25216
rect 14577 25182 14631 25216
rect 13951 25126 14631 25182
rect 13951 25092 14003 25126
rect 14037 25092 14093 25126
rect 14127 25092 14183 25126
rect 14217 25092 14273 25126
rect 14307 25092 14363 25126
rect 14397 25092 14453 25126
rect 14487 25092 14543 25126
rect 14577 25092 14631 25126
rect 13951 25036 14631 25092
rect 13951 25002 14003 25036
rect 14037 25002 14093 25036
rect 14127 25002 14183 25036
rect 14217 25002 14273 25036
rect 14307 25002 14363 25036
rect 14397 25002 14453 25036
rect 14487 25002 14543 25036
rect 14577 25002 14631 25036
rect 13951 24946 14631 25002
rect 13951 24912 14003 24946
rect 14037 24912 14093 24946
rect 14127 24912 14183 24946
rect 14217 24912 14273 24946
rect 14307 24912 14363 24946
rect 14397 24912 14453 24946
rect 14487 24912 14543 24946
rect 14577 24912 14631 24946
rect 13951 24856 14631 24912
rect 13951 24822 14003 24856
rect 14037 24822 14093 24856
rect 14127 24822 14183 24856
rect 14217 24822 14273 24856
rect 14307 24822 14363 24856
rect 14397 24822 14453 24856
rect 14487 24822 14543 24856
rect 14577 24822 14631 24856
rect 13951 24766 14631 24822
rect 13951 24732 14003 24766
rect 14037 24732 14093 24766
rect 14127 24732 14183 24766
rect 14217 24732 14273 24766
rect 14307 24732 14363 24766
rect 14397 24732 14453 24766
rect 14487 24732 14543 24766
rect 14577 24732 14631 24766
rect 13951 24676 14631 24732
rect 13951 24642 14003 24676
rect 14037 24642 14093 24676
rect 14127 24642 14183 24676
rect 14217 24642 14273 24676
rect 14307 24642 14363 24676
rect 14397 24642 14453 24676
rect 14487 24642 14543 24676
rect 14577 24642 14631 24676
rect 13951 24590 14631 24642
rect 15295 25216 15975 25270
rect 15295 25182 15347 25216
rect 15381 25182 15437 25216
rect 15471 25182 15527 25216
rect 15561 25182 15617 25216
rect 15651 25182 15707 25216
rect 15741 25182 15797 25216
rect 15831 25182 15887 25216
rect 15921 25182 15975 25216
rect 15295 25126 15975 25182
rect 15295 25092 15347 25126
rect 15381 25092 15437 25126
rect 15471 25092 15527 25126
rect 15561 25092 15617 25126
rect 15651 25092 15707 25126
rect 15741 25092 15797 25126
rect 15831 25092 15887 25126
rect 15921 25092 15975 25126
rect 15295 25036 15975 25092
rect 15295 25002 15347 25036
rect 15381 25002 15437 25036
rect 15471 25002 15527 25036
rect 15561 25002 15617 25036
rect 15651 25002 15707 25036
rect 15741 25002 15797 25036
rect 15831 25002 15887 25036
rect 15921 25002 15975 25036
rect 15295 24946 15975 25002
rect 15295 24912 15347 24946
rect 15381 24912 15437 24946
rect 15471 24912 15527 24946
rect 15561 24912 15617 24946
rect 15651 24912 15707 24946
rect 15741 24912 15797 24946
rect 15831 24912 15887 24946
rect 15921 24912 15975 24946
rect 15295 24856 15975 24912
rect 15295 24822 15347 24856
rect 15381 24822 15437 24856
rect 15471 24822 15527 24856
rect 15561 24822 15617 24856
rect 15651 24822 15707 24856
rect 15741 24822 15797 24856
rect 15831 24822 15887 24856
rect 15921 24822 15975 24856
rect 15295 24766 15975 24822
rect 15295 24732 15347 24766
rect 15381 24732 15437 24766
rect 15471 24732 15527 24766
rect 15561 24732 15617 24766
rect 15651 24732 15707 24766
rect 15741 24732 15797 24766
rect 15831 24732 15887 24766
rect 15921 24732 15975 24766
rect 15295 24676 15975 24732
rect 15295 24642 15347 24676
rect 15381 24642 15437 24676
rect 15471 24642 15527 24676
rect 15561 24642 15617 24676
rect 15651 24642 15707 24676
rect 15741 24642 15797 24676
rect 15831 24642 15887 24676
rect 15921 24642 15975 24676
rect 15295 24590 15975 24642
rect 16639 25216 17319 25270
rect 16639 25182 16691 25216
rect 16725 25182 16781 25216
rect 16815 25182 16871 25216
rect 16905 25182 16961 25216
rect 16995 25182 17051 25216
rect 17085 25182 17141 25216
rect 17175 25182 17231 25216
rect 17265 25182 17319 25216
rect 16639 25126 17319 25182
rect 16639 25092 16691 25126
rect 16725 25092 16781 25126
rect 16815 25092 16871 25126
rect 16905 25092 16961 25126
rect 16995 25092 17051 25126
rect 17085 25092 17141 25126
rect 17175 25092 17231 25126
rect 17265 25092 17319 25126
rect 16639 25036 17319 25092
rect 16639 25002 16691 25036
rect 16725 25002 16781 25036
rect 16815 25002 16871 25036
rect 16905 25002 16961 25036
rect 16995 25002 17051 25036
rect 17085 25002 17141 25036
rect 17175 25002 17231 25036
rect 17265 25002 17319 25036
rect 16639 24946 17319 25002
rect 16639 24912 16691 24946
rect 16725 24912 16781 24946
rect 16815 24912 16871 24946
rect 16905 24912 16961 24946
rect 16995 24912 17051 24946
rect 17085 24912 17141 24946
rect 17175 24912 17231 24946
rect 17265 24912 17319 24946
rect 16639 24856 17319 24912
rect 16639 24822 16691 24856
rect 16725 24822 16781 24856
rect 16815 24822 16871 24856
rect 16905 24822 16961 24856
rect 16995 24822 17051 24856
rect 17085 24822 17141 24856
rect 17175 24822 17231 24856
rect 17265 24822 17319 24856
rect 16639 24766 17319 24822
rect 16639 24732 16691 24766
rect 16725 24732 16781 24766
rect 16815 24732 16871 24766
rect 16905 24732 16961 24766
rect 16995 24732 17051 24766
rect 17085 24732 17141 24766
rect 17175 24732 17231 24766
rect 17265 24732 17319 24766
rect 16639 24676 17319 24732
rect 16639 24642 16691 24676
rect 16725 24642 16781 24676
rect 16815 24642 16871 24676
rect 16905 24642 16961 24676
rect 16995 24642 17051 24676
rect 17085 24642 17141 24676
rect 17175 24642 17231 24676
rect 17265 24642 17319 24676
rect 16639 24590 17319 24642
<< mvndiff >>
rect 6152 24102 6252 24114
rect 6152 24068 6164 24102
rect 6240 24068 6252 24102
rect 6152 24056 6252 24068
rect 6152 20044 6252 20056
rect 6152 20010 6164 20044
rect 6240 20010 6252 20044
rect 6152 19998 6252 20010
rect 6638 24102 6738 24114
rect 6638 24068 6650 24102
rect 6726 24068 6738 24102
rect 6638 24056 6738 24068
rect 6638 20044 6738 20056
rect 6638 20010 6650 20044
rect 6726 20010 6738 20044
rect 6638 19998 6738 20010
rect 7124 24102 7224 24114
rect 7124 24068 7136 24102
rect 7212 24068 7224 24102
rect 7124 24056 7224 24068
rect 7124 20044 7224 20056
rect 7124 20010 7136 20044
rect 7212 20010 7224 20044
rect 7124 19998 7224 20010
rect 7610 24102 7710 24114
rect 7610 24068 7622 24102
rect 7698 24068 7710 24102
rect 7610 24056 7710 24068
rect 7610 20044 7710 20056
rect 7610 20010 7622 20044
rect 7698 20010 7710 20044
rect 7610 19998 7710 20010
rect 8096 24102 8196 24114
rect 8096 24068 8108 24102
rect 8184 24068 8196 24102
rect 8096 24056 8196 24068
rect 8096 20044 8196 20056
rect 8096 20010 8108 20044
rect 8184 20010 8196 20044
rect 8096 19998 8196 20010
rect 8582 24102 8682 24114
rect 8582 24068 8594 24102
rect 8670 24068 8682 24102
rect 8582 24056 8682 24068
rect 8582 20044 8682 20056
rect 8582 20010 8594 20044
rect 8670 20010 8682 20044
rect 8582 19998 8682 20010
rect 9068 24102 9168 24114
rect 9068 24068 9080 24102
rect 9156 24068 9168 24102
rect 9068 24056 9168 24068
rect 9068 20044 9168 20056
rect 9068 20010 9080 20044
rect 9156 20010 9168 20044
rect 9068 19998 9168 20010
rect 9554 24102 9654 24114
rect 9554 24068 9566 24102
rect 9642 24068 9654 24102
rect 9554 24056 9654 24068
rect 9554 20044 9654 20056
rect 9554 20010 9566 20044
rect 9642 20010 9654 20044
rect 9554 19998 9654 20010
rect 10040 24102 10140 24114
rect 10040 24068 10052 24102
rect 10128 24068 10140 24102
rect 10040 24056 10140 24068
rect 10040 20044 10140 20056
rect 10040 20010 10052 20044
rect 10128 20010 10140 20044
rect 10040 19998 10140 20010
rect 10526 24102 10626 24114
rect 10526 24068 10538 24102
rect 10614 24068 10626 24102
rect 10526 24056 10626 24068
rect 10526 20044 10626 20056
rect 10526 20010 10538 20044
rect 10614 20010 10626 20044
rect 10526 19998 10626 20010
rect 11329 23207 11387 23219
rect 11329 22631 11341 23207
rect 11375 22631 11387 23207
rect 11329 22619 11387 22631
rect 15387 23207 15445 23219
rect 15387 22631 15399 23207
rect 15433 22631 15445 23207
rect 15387 22619 15445 22631
rect 15785 23607 15843 23619
rect 15785 22631 15797 23607
rect 15831 22631 15843 23607
rect 15785 22619 15843 22631
rect 19843 23607 19901 23619
rect 19843 22631 19855 23607
rect 19889 22631 19901 23607
rect 19843 22619 19901 22631
rect 11336 21935 11394 21947
rect 11336 20959 11348 21935
rect 11382 20959 11394 21935
rect 11336 20947 11394 20959
rect 15394 21935 15452 21947
rect 15394 20959 15406 21935
rect 15440 20959 15452 21935
rect 15394 20947 15452 20959
rect 15785 21935 15843 21947
rect 15785 21359 15797 21935
rect 15831 21359 15843 21935
rect 15785 21347 15843 21359
rect 19843 21935 19901 21947
rect 19843 21359 19855 21935
rect 19889 21359 19901 21935
rect 19843 21347 19901 21359
rect 11405 9638 11463 9650
rect 11405 9462 11417 9638
rect 11451 9462 11463 9638
rect 11405 9450 11463 9462
rect 11563 9638 11621 9650
rect 11563 9462 11575 9638
rect 11609 9462 11621 9638
rect 11563 9450 11621 9462
rect 11961 9638 12019 9650
rect 11961 9462 11973 9638
rect 12007 9462 12019 9638
rect 11961 9450 12019 9462
rect 12119 9638 12177 9650
rect 12119 9462 12131 9638
rect 12165 9462 12177 9638
rect 12119 9450 12177 9462
rect 12517 9638 12575 9650
rect 12517 9462 12529 9638
rect 12563 9462 12575 9638
rect 12517 9450 12575 9462
rect 12675 9638 12733 9650
rect 12675 9462 12687 9638
rect 12721 9462 12733 9638
rect 12675 9450 12733 9462
rect 13073 9638 13131 9650
rect 13073 9462 13085 9638
rect 13119 9462 13131 9638
rect 13073 9450 13131 9462
rect 13231 9638 13289 9650
rect 13231 9462 13243 9638
rect 13277 9462 13289 9638
rect 13231 9450 13289 9462
rect 5453 8387 5511 8399
rect 5453 8211 5465 8387
rect 5499 8211 5511 8387
rect 5453 8199 5511 8211
rect 6711 8387 6769 8399
rect 6711 8211 6723 8387
rect 6757 8211 6769 8387
rect 6711 8199 6769 8211
rect 7109 8387 7167 8399
rect 7109 8211 7121 8387
rect 7155 8211 7167 8387
rect 7109 8199 7167 8211
rect 8367 8387 8425 8399
rect 8367 8211 8379 8387
rect 8413 8211 8425 8387
rect 8367 8199 8425 8211
rect 9039 8387 9097 8399
rect 9039 8211 9051 8387
rect 9085 8211 9097 8387
rect 9039 8199 9097 8211
rect 9537 8387 9595 8399
rect 9537 8211 9549 8387
rect 9583 8211 9595 8387
rect 9537 8199 9595 8211
rect 10011 8388 10069 8400
rect 10011 8212 10023 8388
rect 10057 8212 10069 8388
rect 10011 8200 10069 8212
rect 10509 8388 10567 8400
rect 10509 8212 10521 8388
rect 10555 8212 10567 8388
rect 10509 8200 10567 8212
rect 5453 7671 5511 7683
rect 5453 7495 5465 7671
rect 5499 7495 5511 7671
rect 5453 7483 5511 7495
rect 6711 7671 6769 7683
rect 6711 7495 6723 7671
rect 6757 7495 6769 7671
rect 6711 7483 6769 7495
rect 7109 7671 7167 7683
rect 7109 7495 7121 7671
rect 7155 7495 7167 7671
rect 7109 7483 7167 7495
rect 8367 7671 8425 7683
rect 8367 7495 8379 7671
rect 8413 7495 8425 7671
rect 8367 7483 8425 7495
rect 5453 6955 5511 6967
rect 5453 6779 5465 6955
rect 5499 6779 5511 6955
rect 5453 6767 5511 6779
rect 6711 6955 6769 6967
rect 6711 6779 6723 6955
rect 6757 6779 6769 6955
rect 6711 6767 6769 6779
rect 7109 6955 7167 6967
rect 7109 6779 7121 6955
rect 7155 6779 7167 6955
rect 7109 6767 7167 6779
rect 8367 6955 8425 6967
rect 8367 6779 8379 6955
rect 8413 6779 8425 6955
rect 8367 6767 8425 6779
rect 16597 9676 16655 9688
rect 16597 7700 16609 9676
rect 16643 7700 16655 9676
rect 16597 7688 16655 7700
rect 16755 9676 16813 9688
rect 16755 7700 16767 9676
rect 16801 7700 16813 9676
rect 16755 7688 16813 7700
rect 16913 9676 16971 9688
rect 16913 7700 16925 9676
rect 16959 7700 16971 9676
rect 16913 7688 16971 7700
rect 17071 9676 17129 9688
rect 17071 7700 17083 9676
rect 17117 7700 17129 9676
rect 17071 7688 17129 7700
rect 17229 9676 17287 9688
rect 17229 7700 17241 9676
rect 17275 7700 17287 9676
rect 17229 7688 17287 7700
rect 17387 9676 17445 9688
rect 17387 7700 17399 9676
rect 17433 7700 17445 9676
rect 17387 7688 17445 7700
rect 17545 9676 17603 9688
rect 17545 7700 17557 9676
rect 17591 7700 17603 9676
rect 17545 7688 17603 7700
rect 17703 9676 17761 9688
rect 17703 7700 17715 9676
rect 17749 7700 17761 9676
rect 17703 7688 17761 7700
rect 17861 9676 17919 9688
rect 17861 7700 17873 9676
rect 17907 7700 17919 9676
rect 17861 7688 17919 7700
rect 18019 9676 18077 9688
rect 18019 7700 18031 9676
rect 18065 7700 18077 9676
rect 18019 7688 18077 7700
rect 18177 9676 18235 9688
rect 18177 7700 18189 9676
rect 18223 7700 18235 9676
rect 18177 7688 18235 7700
rect 18335 9676 18393 9688
rect 18335 7700 18347 9676
rect 18381 7700 18393 9676
rect 18335 7688 18393 7700
rect 18493 9676 18551 9688
rect 18493 7700 18505 9676
rect 18539 7700 18551 9676
rect 18493 7688 18551 7700
rect 18651 9676 18709 9688
rect 18651 7700 18663 9676
rect 18697 7700 18709 9676
rect 18651 7688 18709 7700
rect 18809 9676 18867 9688
rect 18809 7700 18821 9676
rect 18855 7700 18867 9676
rect 18809 7688 18867 7700
rect 18967 9676 19025 9688
rect 18967 7700 18979 9676
rect 19013 7700 19025 9676
rect 18967 7688 19025 7700
rect 19125 9676 19183 9688
rect 19125 7700 19137 9676
rect 19171 7700 19183 9676
rect 19125 7688 19183 7700
rect 19283 9676 19341 9688
rect 19283 7700 19295 9676
rect 19329 7700 19341 9676
rect 19283 7688 19341 7700
rect 19441 9676 19499 9688
rect 19441 7700 19453 9676
rect 19487 7700 19499 9676
rect 19441 7688 19499 7700
rect 19599 9676 19657 9688
rect 19599 7700 19611 9676
rect 19645 7700 19657 9676
rect 19599 7688 19657 7700
rect 19757 9676 19815 9688
rect 19757 7700 19769 9676
rect 19803 7700 19815 9676
rect 19757 7688 19815 7700
rect 19915 9676 19973 9688
rect 19915 7700 19927 9676
rect 19961 7700 19973 9676
rect 19915 7688 19973 7700
rect 20073 9676 20131 9688
rect 20073 7700 20085 9676
rect 20119 7700 20131 9676
rect 20073 7688 20131 7700
rect 5453 6239 5511 6251
rect 5453 6063 5465 6239
rect 5499 6063 5511 6239
rect 5453 6051 5511 6063
rect 6711 6239 6769 6251
rect 6711 6063 6723 6239
rect 6757 6063 6769 6239
rect 6711 6051 6769 6063
rect 7109 6239 7167 6251
rect 7109 6063 7121 6239
rect 7155 6063 7167 6239
rect 7109 6051 7167 6063
rect 8367 6239 8425 6251
rect 8367 6063 8379 6239
rect 8413 6063 8425 6239
rect 8367 6051 8425 6063
rect 16681 7177 16881 7189
rect 16681 7143 16693 7177
rect 16869 7143 16881 7177
rect 16681 7131 16881 7143
rect 16681 5119 16881 5131
rect 16681 5085 16693 5119
rect 16869 5085 16881 5119
rect 16681 5073 16881 5085
rect 17267 7177 17467 7189
rect 17267 7143 17279 7177
rect 17455 7143 17467 7177
rect 17267 7131 17467 7143
rect 17267 5119 17467 5131
rect 17267 5085 17279 5119
rect 17455 5085 17467 5119
rect 17267 5073 17467 5085
rect 17853 7177 18053 7189
rect 17853 7143 17865 7177
rect 18041 7143 18053 7177
rect 17853 7131 18053 7143
rect 17853 5119 18053 5131
rect 17853 5085 17865 5119
rect 18041 5085 18053 5119
rect 17853 5073 18053 5085
rect 16681 4715 16881 4727
rect 16681 4681 16693 4715
rect 16869 4681 16881 4715
rect 16681 4669 16881 4681
rect 16681 2657 16881 2669
rect 16681 2623 16693 2657
rect 16869 2623 16881 2657
rect 16681 2611 16881 2623
rect 17267 4715 17467 4727
rect 17267 4681 17279 4715
rect 17455 4681 17467 4715
rect 17267 4669 17467 4681
rect 17267 2657 17467 2669
rect 17267 2623 17279 2657
rect 17455 2623 17467 2657
rect 17267 2611 17467 2623
rect 17853 4715 18053 4727
rect 17853 4681 17865 4715
rect 18041 4681 18053 4715
rect 17853 4669 18053 4681
rect 17853 2657 18053 2669
rect 17853 2623 17865 2657
rect 18041 2623 18053 2657
rect 17853 2611 18053 2623
rect 21737 7945 23737 7957
rect 21737 7911 21749 7945
rect 23725 7911 23737 7945
rect 21737 7899 23737 7911
rect 21737 6087 23737 6099
rect 21737 6053 21749 6087
rect 23725 6053 23737 6087
rect 21737 6041 23737 6053
rect 21737 5695 23737 5707
rect 21737 5661 21749 5695
rect 23725 5661 23737 5695
rect 21737 5649 23737 5661
rect 21737 3837 23737 3849
rect 21737 3803 21749 3837
rect 23725 3803 23737 3837
rect 21737 3791 23737 3803
rect 21434 2915 21492 2927
rect 21434 1939 21446 2915
rect 21480 1939 21492 2915
rect 21434 1927 21492 1939
rect 21692 2915 21750 2927
rect 21692 1939 21704 2915
rect 21738 1939 21750 2915
rect 21692 1927 21750 1939
rect 21950 2915 22008 2927
rect 21950 1939 21962 2915
rect 21996 1939 22008 2915
rect 21950 1927 22008 1939
rect 22208 2915 22266 2927
rect 22208 1939 22220 2915
rect 22254 1939 22266 2915
rect 22208 1927 22266 1939
rect 22466 2915 22524 2927
rect 22466 1939 22478 2915
rect 22512 1939 22524 2915
rect 22466 1927 22524 1939
rect 22724 2915 22782 2927
rect 22724 1939 22736 2915
rect 22770 1939 22782 2915
rect 22724 1927 22782 1939
rect 22982 2915 23040 2927
rect 22982 1939 22994 2915
rect 23028 1939 23040 2915
rect 22982 1927 23040 1939
rect 23240 2915 23298 2927
rect 23240 1939 23252 2915
rect 23286 1939 23298 2915
rect 23240 1927 23298 1939
rect 23498 2915 23556 2927
rect 23498 1939 23510 2915
rect 23544 1939 23556 2915
rect 23498 1927 23556 1939
rect 23756 2915 23814 2927
rect 23756 1939 23768 2915
rect 23802 1939 23814 2915
rect 23756 1927 23814 1939
rect 24014 2915 24072 2927
rect 24014 1939 24026 2915
rect 24060 1939 24072 2915
rect 24014 1927 24072 1939
rect 24666 3837 26666 3849
rect 24666 3803 24678 3837
rect 26654 3803 26666 3837
rect 24666 3791 26666 3803
rect 24666 1979 26666 1991
rect 24666 1945 24678 1979
rect 26654 1945 26666 1979
rect 24666 1933 26666 1945
<< mvpdiff >>
rect 6221 30906 6279 30918
rect 6221 30730 6233 30906
rect 6267 30730 6279 30906
rect 6221 30718 6279 30730
rect 8279 30906 8337 30918
rect 8279 30730 8291 30906
rect 8325 30730 8337 30906
rect 8279 30718 8337 30730
rect 8547 30906 8605 30918
rect 8547 30730 8559 30906
rect 8593 30730 8605 30906
rect 8547 30718 8605 30730
rect 10605 30906 10663 30918
rect 10605 30730 10617 30906
rect 10651 30730 10663 30906
rect 10605 30718 10663 30730
rect 6346 19039 6404 19051
rect 6346 18763 6358 19039
rect 6392 18763 6404 19039
rect 6346 18751 6404 18763
rect 10404 19039 10462 19051
rect 10404 18763 10416 19039
rect 10450 18763 10462 19039
rect 10404 18751 10462 18763
rect 6346 18503 6404 18515
rect 6346 18227 6358 18503
rect 6392 18227 6404 18503
rect 6346 18215 6404 18227
rect 10404 18503 10462 18515
rect 10404 18227 10416 18503
rect 10450 18227 10462 18503
rect 10404 18215 10462 18227
rect 6346 17639 6404 17651
rect 6346 17063 6358 17639
rect 6392 17063 6404 17639
rect 6346 17051 6404 17063
rect 10404 17639 10462 17651
rect 10404 17063 10416 17639
rect 10450 17063 10462 17639
rect 10404 17051 10462 17063
rect 11434 19039 11492 19051
rect 11434 17063 11446 19039
rect 11480 17063 11492 19039
rect 11434 17051 11492 17063
rect 15492 19039 15550 19051
rect 15492 17063 15504 19039
rect 15538 17063 15550 19039
rect 15492 17051 15550 17063
rect 15760 19039 15818 19051
rect 15760 17063 15772 19039
rect 15806 17063 15818 19039
rect 15760 17051 15818 17063
rect 19818 19039 19876 19051
rect 19818 17063 19830 19039
rect 19864 17063 19876 19039
rect 19818 17051 19876 17063
rect 8356 14835 8414 14847
rect 8356 14659 8368 14835
rect 8402 14659 8414 14835
rect 8356 14647 8414 14659
rect 10404 14835 10462 14847
rect 10404 14659 10416 14835
rect 10450 14659 10462 14835
rect 10404 14647 10462 14659
rect 11434 16635 11492 16647
rect 11434 14659 11446 16635
rect 11480 14659 11492 16635
rect 11434 14647 11492 14659
rect 15492 16635 15550 16647
rect 15492 14659 15504 16635
rect 15538 14659 15550 16635
rect 15492 14647 15550 14659
rect 15760 16635 15818 16647
rect 15760 14659 15772 16635
rect 15806 14659 15818 16635
rect 15760 14647 15818 14659
rect 19818 16635 19876 16647
rect 19818 14659 19830 16635
rect 19864 14659 19876 16635
rect 19818 14647 19876 14659
rect 20899 18768 20999 18780
rect 20899 18734 20911 18768
rect 20987 18734 20999 18768
rect 20899 18722 20999 18734
rect 20899 14710 20999 14722
rect 20899 14676 20911 14710
rect 20987 14676 20999 14710
rect 20899 14664 20999 14676
rect 21403 18768 21503 18780
rect 21403 18734 21415 18768
rect 21491 18734 21503 18768
rect 21403 18722 21503 18734
rect 21403 14710 21503 14722
rect 21403 14676 21415 14710
rect 21491 14676 21503 14710
rect 21403 14664 21503 14676
rect 8061 12311 8119 12323
rect 8061 12135 8073 12311
rect 8107 12135 8119 12311
rect 8061 12123 8119 12135
rect 10129 12311 10187 12323
rect 10129 12135 10141 12311
rect 10175 12135 10187 12311
rect 10129 12123 10187 12135
rect 6061 11548 6119 11560
rect 6061 11172 6073 11548
rect 6107 11172 6119 11548
rect 6061 11160 6119 11172
rect 10119 11548 10177 11560
rect 10119 11172 10131 11548
rect 10165 11172 10177 11548
rect 10119 11160 10177 11172
rect 6173 10562 6231 10574
rect 6173 10086 6185 10562
rect 6219 10086 6231 10562
rect 6173 10074 6231 10086
rect 6711 10562 6769 10574
rect 6711 10086 6723 10562
rect 6757 10086 6769 10562
rect 6711 10074 6769 10086
rect 7109 10562 7167 10574
rect 7109 10086 7121 10562
rect 7155 10086 7167 10562
rect 7109 10074 7167 10086
rect 7647 10562 7705 10574
rect 7647 10086 7659 10562
rect 7693 10086 7705 10562
rect 7647 10074 7705 10086
rect 9039 10580 9097 10592
rect 9039 10104 9051 10580
rect 9085 10104 9097 10580
rect 9039 10092 9097 10104
rect 9577 10580 9635 10592
rect 9577 10104 9589 10580
rect 9623 10104 9635 10580
rect 9577 10092 9635 10104
rect 9971 10580 10029 10592
rect 9971 10104 9983 10580
rect 10017 10104 10029 10580
rect 9971 10092 10029 10104
rect 10509 10580 10567 10592
rect 10509 10104 10521 10580
rect 10555 10104 10567 10580
rect 10509 10092 10567 10104
rect 12021 10853 12079 10865
rect 12021 10677 12033 10853
rect 12067 10677 12079 10853
rect 12021 10665 12079 10677
rect 12179 10853 12237 10865
rect 12179 10677 12191 10853
rect 12225 10677 12237 10853
rect 12179 10665 12237 10677
rect 12337 10853 12395 10865
rect 12337 10677 12349 10853
rect 12383 10677 12395 10853
rect 12337 10665 12395 10677
rect 12495 10853 12553 10865
rect 12495 10677 12507 10853
rect 12541 10677 12553 10853
rect 12495 10665 12553 10677
rect 12653 10853 12711 10865
rect 12653 10677 12665 10853
rect 12699 10677 12711 10853
rect 12653 10665 12711 10677
rect 6173 9520 6231 9532
rect 6173 9044 6185 9520
rect 6219 9044 6231 9520
rect 6173 9032 6231 9044
rect 6711 9520 6769 9532
rect 6711 9044 6723 9520
rect 6757 9044 6769 9520
rect 6711 9032 6769 9044
rect 7109 9520 7167 9532
rect 7109 9044 7121 9520
rect 7155 9044 7167 9520
rect 7109 9032 7167 9044
rect 7647 9520 7705 9532
rect 7647 9044 7659 9520
rect 7693 9044 7705 9520
rect 7647 9032 7705 9044
rect 9039 9495 9097 9507
rect 9039 9019 9051 9495
rect 9085 9019 9097 9495
rect 9039 9007 9097 9019
rect 9577 9495 9635 9507
rect 9577 9019 9589 9495
rect 9623 9019 9635 9495
rect 9577 9007 9635 9019
rect 9971 9495 10029 9507
rect 9971 9019 9983 9495
rect 10017 9019 10029 9495
rect 9971 9007 10029 9019
rect 10509 9495 10567 9507
rect 10509 9019 10521 9495
rect 10555 9019 10567 9495
rect 10509 9007 10567 9019
rect 24831 7945 25631 7957
rect 24831 7911 24843 7945
rect 25619 7911 25631 7945
rect 24831 7899 25631 7911
rect 24831 7687 25631 7699
rect 24831 7653 24843 7687
rect 25619 7653 25631 7687
rect 24831 7641 25631 7653
rect 24831 7239 26531 7251
rect 24831 7205 24843 7239
rect 26519 7205 26531 7239
rect 24831 7193 26531 7205
rect 24831 6981 26531 6993
rect 24831 6947 24843 6981
rect 26519 6947 26531 6981
rect 24831 6935 26531 6947
rect 24831 6723 26531 6735
rect 24831 6689 24843 6723
rect 26519 6689 26531 6723
rect 24831 6677 26531 6689
rect 24831 6465 26531 6477
rect 24831 6431 24843 6465
rect 26519 6431 26531 6465
rect 24831 6419 26531 6431
rect 24831 6207 26531 6219
rect 24831 6173 24843 6207
rect 26519 6173 26531 6207
rect 24831 6161 26531 6173
rect 24831 5949 26531 5961
rect 24831 5915 24843 5949
rect 26519 5915 26531 5949
rect 24831 5903 26531 5915
rect 24831 5691 26531 5703
rect 24831 5657 24843 5691
rect 26519 5657 26531 5691
rect 24831 5645 26531 5657
rect 24831 5433 26531 5445
rect 24831 5399 24843 5433
rect 26519 5399 26531 5433
rect 24831 5387 26531 5399
rect 24831 5175 26531 5187
rect 24831 5141 24843 5175
rect 26519 5141 26531 5175
rect 24831 5129 26531 5141
<< pdiffc >>
rect 14003 27870 14037 27904
rect 14093 27870 14127 27904
rect 14183 27870 14217 27904
rect 14273 27870 14307 27904
rect 14363 27870 14397 27904
rect 14453 27870 14487 27904
rect 14543 27870 14577 27904
rect 14003 27780 14037 27814
rect 14093 27780 14127 27814
rect 14183 27780 14217 27814
rect 14273 27780 14307 27814
rect 14363 27780 14397 27814
rect 14453 27780 14487 27814
rect 14543 27780 14577 27814
rect 14003 27690 14037 27724
rect 14093 27690 14127 27724
rect 14183 27690 14217 27724
rect 14273 27690 14307 27724
rect 14363 27690 14397 27724
rect 14453 27690 14487 27724
rect 14543 27690 14577 27724
rect 14003 27600 14037 27634
rect 14093 27600 14127 27634
rect 14183 27600 14217 27634
rect 14273 27600 14307 27634
rect 14363 27600 14397 27634
rect 14453 27600 14487 27634
rect 14543 27600 14577 27634
rect 14003 27510 14037 27544
rect 14093 27510 14127 27544
rect 14183 27510 14217 27544
rect 14273 27510 14307 27544
rect 14363 27510 14397 27544
rect 14453 27510 14487 27544
rect 14543 27510 14577 27544
rect 14003 27420 14037 27454
rect 14093 27420 14127 27454
rect 14183 27420 14217 27454
rect 14273 27420 14307 27454
rect 14363 27420 14397 27454
rect 14453 27420 14487 27454
rect 14543 27420 14577 27454
rect 14003 27330 14037 27364
rect 14093 27330 14127 27364
rect 14183 27330 14217 27364
rect 14273 27330 14307 27364
rect 14363 27330 14397 27364
rect 14453 27330 14487 27364
rect 14543 27330 14577 27364
rect 15347 27870 15381 27904
rect 15437 27870 15471 27904
rect 15527 27870 15561 27904
rect 15617 27870 15651 27904
rect 15707 27870 15741 27904
rect 15797 27870 15831 27904
rect 15887 27870 15921 27904
rect 15347 27780 15381 27814
rect 15437 27780 15471 27814
rect 15527 27780 15561 27814
rect 15617 27780 15651 27814
rect 15707 27780 15741 27814
rect 15797 27780 15831 27814
rect 15887 27780 15921 27814
rect 15347 27690 15381 27724
rect 15437 27690 15471 27724
rect 15527 27690 15561 27724
rect 15617 27690 15651 27724
rect 15707 27690 15741 27724
rect 15797 27690 15831 27724
rect 15887 27690 15921 27724
rect 15347 27600 15381 27634
rect 15437 27600 15471 27634
rect 15527 27600 15561 27634
rect 15617 27600 15651 27634
rect 15707 27600 15741 27634
rect 15797 27600 15831 27634
rect 15887 27600 15921 27634
rect 15347 27510 15381 27544
rect 15437 27510 15471 27544
rect 15527 27510 15561 27544
rect 15617 27510 15651 27544
rect 15707 27510 15741 27544
rect 15797 27510 15831 27544
rect 15887 27510 15921 27544
rect 15347 27420 15381 27454
rect 15437 27420 15471 27454
rect 15527 27420 15561 27454
rect 15617 27420 15651 27454
rect 15707 27420 15741 27454
rect 15797 27420 15831 27454
rect 15887 27420 15921 27454
rect 15347 27330 15381 27364
rect 15437 27330 15471 27364
rect 15527 27330 15561 27364
rect 15617 27330 15651 27364
rect 15707 27330 15741 27364
rect 15797 27330 15831 27364
rect 15887 27330 15921 27364
rect 16691 27870 16725 27904
rect 16781 27870 16815 27904
rect 16871 27870 16905 27904
rect 16961 27870 16995 27904
rect 17051 27870 17085 27904
rect 17141 27870 17175 27904
rect 17231 27870 17265 27904
rect 16691 27780 16725 27814
rect 16781 27780 16815 27814
rect 16871 27780 16905 27814
rect 16961 27780 16995 27814
rect 17051 27780 17085 27814
rect 17141 27780 17175 27814
rect 17231 27780 17265 27814
rect 16691 27690 16725 27724
rect 16781 27690 16815 27724
rect 16871 27690 16905 27724
rect 16961 27690 16995 27724
rect 17051 27690 17085 27724
rect 17141 27690 17175 27724
rect 17231 27690 17265 27724
rect 16691 27600 16725 27634
rect 16781 27600 16815 27634
rect 16871 27600 16905 27634
rect 16961 27600 16995 27634
rect 17051 27600 17085 27634
rect 17141 27600 17175 27634
rect 17231 27600 17265 27634
rect 16691 27510 16725 27544
rect 16781 27510 16815 27544
rect 16871 27510 16905 27544
rect 16961 27510 16995 27544
rect 17051 27510 17085 27544
rect 17141 27510 17175 27544
rect 17231 27510 17265 27544
rect 16691 27420 16725 27454
rect 16781 27420 16815 27454
rect 16871 27420 16905 27454
rect 16961 27420 16995 27454
rect 17051 27420 17085 27454
rect 17141 27420 17175 27454
rect 17231 27420 17265 27454
rect 16691 27330 16725 27364
rect 16781 27330 16815 27364
rect 16871 27330 16905 27364
rect 16961 27330 16995 27364
rect 17051 27330 17085 27364
rect 17141 27330 17175 27364
rect 17231 27330 17265 27364
rect 14003 26526 14037 26560
rect 14093 26526 14127 26560
rect 14183 26526 14217 26560
rect 14273 26526 14307 26560
rect 14363 26526 14397 26560
rect 14453 26526 14487 26560
rect 14543 26526 14577 26560
rect 14003 26436 14037 26470
rect 14093 26436 14127 26470
rect 14183 26436 14217 26470
rect 14273 26436 14307 26470
rect 14363 26436 14397 26470
rect 14453 26436 14487 26470
rect 14543 26436 14577 26470
rect 14003 26346 14037 26380
rect 14093 26346 14127 26380
rect 14183 26346 14217 26380
rect 14273 26346 14307 26380
rect 14363 26346 14397 26380
rect 14453 26346 14487 26380
rect 14543 26346 14577 26380
rect 14003 26256 14037 26290
rect 14093 26256 14127 26290
rect 14183 26256 14217 26290
rect 14273 26256 14307 26290
rect 14363 26256 14397 26290
rect 14453 26256 14487 26290
rect 14543 26256 14577 26290
rect 14003 26166 14037 26200
rect 14093 26166 14127 26200
rect 14183 26166 14217 26200
rect 14273 26166 14307 26200
rect 14363 26166 14397 26200
rect 14453 26166 14487 26200
rect 14543 26166 14577 26200
rect 14003 26076 14037 26110
rect 14093 26076 14127 26110
rect 14183 26076 14217 26110
rect 14273 26076 14307 26110
rect 14363 26076 14397 26110
rect 14453 26076 14487 26110
rect 14543 26076 14577 26110
rect 14003 25986 14037 26020
rect 14093 25986 14127 26020
rect 14183 25986 14217 26020
rect 14273 25986 14307 26020
rect 14363 25986 14397 26020
rect 14453 25986 14487 26020
rect 14543 25986 14577 26020
rect 15347 26526 15381 26560
rect 15437 26526 15471 26560
rect 15527 26526 15561 26560
rect 15617 26526 15651 26560
rect 15707 26526 15741 26560
rect 15797 26526 15831 26560
rect 15887 26526 15921 26560
rect 15347 26436 15381 26470
rect 15437 26436 15471 26470
rect 15527 26436 15561 26470
rect 15617 26436 15651 26470
rect 15707 26436 15741 26470
rect 15797 26436 15831 26470
rect 15887 26436 15921 26470
rect 15347 26346 15381 26380
rect 15437 26346 15471 26380
rect 15527 26346 15561 26380
rect 15617 26346 15651 26380
rect 15707 26346 15741 26380
rect 15797 26346 15831 26380
rect 15887 26346 15921 26380
rect 15347 26256 15381 26290
rect 15437 26256 15471 26290
rect 15527 26256 15561 26290
rect 15617 26256 15651 26290
rect 15707 26256 15741 26290
rect 15797 26256 15831 26290
rect 15887 26256 15921 26290
rect 15347 26166 15381 26200
rect 15437 26166 15471 26200
rect 15527 26166 15561 26200
rect 15617 26166 15651 26200
rect 15707 26166 15741 26200
rect 15797 26166 15831 26200
rect 15887 26166 15921 26200
rect 15347 26076 15381 26110
rect 15437 26076 15471 26110
rect 15527 26076 15561 26110
rect 15617 26076 15651 26110
rect 15707 26076 15741 26110
rect 15797 26076 15831 26110
rect 15887 26076 15921 26110
rect 15347 25986 15381 26020
rect 15437 25986 15471 26020
rect 15527 25986 15561 26020
rect 15617 25986 15651 26020
rect 15707 25986 15741 26020
rect 15797 25986 15831 26020
rect 15887 25986 15921 26020
rect 16691 26526 16725 26560
rect 16781 26526 16815 26560
rect 16871 26526 16905 26560
rect 16961 26526 16995 26560
rect 17051 26526 17085 26560
rect 17141 26526 17175 26560
rect 17231 26526 17265 26560
rect 16691 26436 16725 26470
rect 16781 26436 16815 26470
rect 16871 26436 16905 26470
rect 16961 26436 16995 26470
rect 17051 26436 17085 26470
rect 17141 26436 17175 26470
rect 17231 26436 17265 26470
rect 16691 26346 16725 26380
rect 16781 26346 16815 26380
rect 16871 26346 16905 26380
rect 16961 26346 16995 26380
rect 17051 26346 17085 26380
rect 17141 26346 17175 26380
rect 17231 26346 17265 26380
rect 16691 26256 16725 26290
rect 16781 26256 16815 26290
rect 16871 26256 16905 26290
rect 16961 26256 16995 26290
rect 17051 26256 17085 26290
rect 17141 26256 17175 26290
rect 17231 26256 17265 26290
rect 16691 26166 16725 26200
rect 16781 26166 16815 26200
rect 16871 26166 16905 26200
rect 16961 26166 16995 26200
rect 17051 26166 17085 26200
rect 17141 26166 17175 26200
rect 17231 26166 17265 26200
rect 16691 26076 16725 26110
rect 16781 26076 16815 26110
rect 16871 26076 16905 26110
rect 16961 26076 16995 26110
rect 17051 26076 17085 26110
rect 17141 26076 17175 26110
rect 17231 26076 17265 26110
rect 16691 25986 16725 26020
rect 16781 25986 16815 26020
rect 16871 25986 16905 26020
rect 16961 25986 16995 26020
rect 17051 25986 17085 26020
rect 17141 25986 17175 26020
rect 17231 25986 17265 26020
rect 14003 25182 14037 25216
rect 14093 25182 14127 25216
rect 14183 25182 14217 25216
rect 14273 25182 14307 25216
rect 14363 25182 14397 25216
rect 14453 25182 14487 25216
rect 14543 25182 14577 25216
rect 14003 25092 14037 25126
rect 14093 25092 14127 25126
rect 14183 25092 14217 25126
rect 14273 25092 14307 25126
rect 14363 25092 14397 25126
rect 14453 25092 14487 25126
rect 14543 25092 14577 25126
rect 14003 25002 14037 25036
rect 14093 25002 14127 25036
rect 14183 25002 14217 25036
rect 14273 25002 14307 25036
rect 14363 25002 14397 25036
rect 14453 25002 14487 25036
rect 14543 25002 14577 25036
rect 14003 24912 14037 24946
rect 14093 24912 14127 24946
rect 14183 24912 14217 24946
rect 14273 24912 14307 24946
rect 14363 24912 14397 24946
rect 14453 24912 14487 24946
rect 14543 24912 14577 24946
rect 14003 24822 14037 24856
rect 14093 24822 14127 24856
rect 14183 24822 14217 24856
rect 14273 24822 14307 24856
rect 14363 24822 14397 24856
rect 14453 24822 14487 24856
rect 14543 24822 14577 24856
rect 14003 24732 14037 24766
rect 14093 24732 14127 24766
rect 14183 24732 14217 24766
rect 14273 24732 14307 24766
rect 14363 24732 14397 24766
rect 14453 24732 14487 24766
rect 14543 24732 14577 24766
rect 14003 24642 14037 24676
rect 14093 24642 14127 24676
rect 14183 24642 14217 24676
rect 14273 24642 14307 24676
rect 14363 24642 14397 24676
rect 14453 24642 14487 24676
rect 14543 24642 14577 24676
rect 15347 25182 15381 25216
rect 15437 25182 15471 25216
rect 15527 25182 15561 25216
rect 15617 25182 15651 25216
rect 15707 25182 15741 25216
rect 15797 25182 15831 25216
rect 15887 25182 15921 25216
rect 15347 25092 15381 25126
rect 15437 25092 15471 25126
rect 15527 25092 15561 25126
rect 15617 25092 15651 25126
rect 15707 25092 15741 25126
rect 15797 25092 15831 25126
rect 15887 25092 15921 25126
rect 15347 25002 15381 25036
rect 15437 25002 15471 25036
rect 15527 25002 15561 25036
rect 15617 25002 15651 25036
rect 15707 25002 15741 25036
rect 15797 25002 15831 25036
rect 15887 25002 15921 25036
rect 15347 24912 15381 24946
rect 15437 24912 15471 24946
rect 15527 24912 15561 24946
rect 15617 24912 15651 24946
rect 15707 24912 15741 24946
rect 15797 24912 15831 24946
rect 15887 24912 15921 24946
rect 15347 24822 15381 24856
rect 15437 24822 15471 24856
rect 15527 24822 15561 24856
rect 15617 24822 15651 24856
rect 15707 24822 15741 24856
rect 15797 24822 15831 24856
rect 15887 24822 15921 24856
rect 15347 24732 15381 24766
rect 15437 24732 15471 24766
rect 15527 24732 15561 24766
rect 15617 24732 15651 24766
rect 15707 24732 15741 24766
rect 15797 24732 15831 24766
rect 15887 24732 15921 24766
rect 15347 24642 15381 24676
rect 15437 24642 15471 24676
rect 15527 24642 15561 24676
rect 15617 24642 15651 24676
rect 15707 24642 15741 24676
rect 15797 24642 15831 24676
rect 15887 24642 15921 24676
rect 16691 25182 16725 25216
rect 16781 25182 16815 25216
rect 16871 25182 16905 25216
rect 16961 25182 16995 25216
rect 17051 25182 17085 25216
rect 17141 25182 17175 25216
rect 17231 25182 17265 25216
rect 16691 25092 16725 25126
rect 16781 25092 16815 25126
rect 16871 25092 16905 25126
rect 16961 25092 16995 25126
rect 17051 25092 17085 25126
rect 17141 25092 17175 25126
rect 17231 25092 17265 25126
rect 16691 25002 16725 25036
rect 16781 25002 16815 25036
rect 16871 25002 16905 25036
rect 16961 25002 16995 25036
rect 17051 25002 17085 25036
rect 17141 25002 17175 25036
rect 17231 25002 17265 25036
rect 16691 24912 16725 24946
rect 16781 24912 16815 24946
rect 16871 24912 16905 24946
rect 16961 24912 16995 24946
rect 17051 24912 17085 24946
rect 17141 24912 17175 24946
rect 17231 24912 17265 24946
rect 16691 24822 16725 24856
rect 16781 24822 16815 24856
rect 16871 24822 16905 24856
rect 16961 24822 16995 24856
rect 17051 24822 17085 24856
rect 17141 24822 17175 24856
rect 17231 24822 17265 24856
rect 16691 24732 16725 24766
rect 16781 24732 16815 24766
rect 16871 24732 16905 24766
rect 16961 24732 16995 24766
rect 17051 24732 17085 24766
rect 17141 24732 17175 24766
rect 17231 24732 17265 24766
rect 16691 24642 16725 24676
rect 16781 24642 16815 24676
rect 16871 24642 16905 24676
rect 16961 24642 16995 24676
rect 17051 24642 17085 24676
rect 17141 24642 17175 24676
rect 17231 24642 17265 24676
<< mvndiffc >>
rect 6164 24068 6240 24102
rect 6164 20010 6240 20044
rect 6650 24068 6726 24102
rect 6650 20010 6726 20044
rect 7136 24068 7212 24102
rect 7136 20010 7212 20044
rect 7622 24068 7698 24102
rect 7622 20010 7698 20044
rect 8108 24068 8184 24102
rect 8108 20010 8184 20044
rect 8594 24068 8670 24102
rect 8594 20010 8670 20044
rect 9080 24068 9156 24102
rect 9080 20010 9156 20044
rect 9566 24068 9642 24102
rect 9566 20010 9642 20044
rect 10052 24068 10128 24102
rect 10052 20010 10128 20044
rect 10538 24068 10614 24102
rect 10538 20010 10614 20044
rect 11341 22631 11375 23207
rect 15399 22631 15433 23207
rect 15797 22631 15831 23607
rect 19855 22631 19889 23607
rect 11348 20959 11382 21935
rect 15406 20959 15440 21935
rect 15797 21359 15831 21935
rect 19855 21359 19889 21935
rect 11417 9462 11451 9638
rect 11575 9462 11609 9638
rect 11973 9462 12007 9638
rect 12131 9462 12165 9638
rect 12529 9462 12563 9638
rect 12687 9462 12721 9638
rect 13085 9462 13119 9638
rect 13243 9462 13277 9638
rect 5465 8211 5499 8387
rect 6723 8211 6757 8387
rect 7121 8211 7155 8387
rect 8379 8211 8413 8387
rect 9051 8211 9085 8387
rect 9549 8211 9583 8387
rect 10023 8212 10057 8388
rect 10521 8212 10555 8388
rect 5465 7495 5499 7671
rect 6723 7495 6757 7671
rect 7121 7495 7155 7671
rect 8379 7495 8413 7671
rect 5465 6779 5499 6955
rect 6723 6779 6757 6955
rect 7121 6779 7155 6955
rect 8379 6779 8413 6955
rect 16609 7700 16643 9676
rect 16767 7700 16801 9676
rect 16925 7700 16959 9676
rect 17083 7700 17117 9676
rect 17241 7700 17275 9676
rect 17399 7700 17433 9676
rect 17557 7700 17591 9676
rect 17715 7700 17749 9676
rect 17873 7700 17907 9676
rect 18031 7700 18065 9676
rect 18189 7700 18223 9676
rect 18347 7700 18381 9676
rect 18505 7700 18539 9676
rect 18663 7700 18697 9676
rect 18821 7700 18855 9676
rect 18979 7700 19013 9676
rect 19137 7700 19171 9676
rect 19295 7700 19329 9676
rect 19453 7700 19487 9676
rect 19611 7700 19645 9676
rect 19769 7700 19803 9676
rect 19927 7700 19961 9676
rect 20085 7700 20119 9676
rect 5465 6063 5499 6239
rect 6723 6063 6757 6239
rect 7121 6063 7155 6239
rect 8379 6063 8413 6239
rect 16693 7143 16869 7177
rect 16693 5085 16869 5119
rect 17279 7143 17455 7177
rect 17279 5085 17455 5119
rect 17865 7143 18041 7177
rect 17865 5085 18041 5119
rect 16693 4681 16869 4715
rect 16693 2623 16869 2657
rect 17279 4681 17455 4715
rect 17279 2623 17455 2657
rect 17865 4681 18041 4715
rect 17865 2623 18041 2657
rect 21749 7911 23725 7945
rect 21749 6053 23725 6087
rect 21749 5661 23725 5695
rect 21749 3803 23725 3837
rect 21446 1939 21480 2915
rect 21704 1939 21738 2915
rect 21962 1939 21996 2915
rect 22220 1939 22254 2915
rect 22478 1939 22512 2915
rect 22736 1939 22770 2915
rect 22994 1939 23028 2915
rect 23252 1939 23286 2915
rect 23510 1939 23544 2915
rect 23768 1939 23802 2915
rect 24026 1939 24060 2915
rect 24678 3803 26654 3837
rect 24678 1945 26654 1979
<< mvpdiffc >>
rect 6233 30730 6267 30906
rect 8291 30730 8325 30906
rect 8559 30730 8593 30906
rect 10617 30730 10651 30906
rect 6358 18763 6392 19039
rect 10416 18763 10450 19039
rect 6358 18227 6392 18503
rect 10416 18227 10450 18503
rect 6358 17063 6392 17639
rect 10416 17063 10450 17639
rect 11446 17063 11480 19039
rect 15504 17063 15538 19039
rect 15772 17063 15806 19039
rect 19830 17063 19864 19039
rect 8368 14659 8402 14835
rect 10416 14659 10450 14835
rect 11446 14659 11480 16635
rect 15504 14659 15538 16635
rect 15772 14659 15806 16635
rect 19830 14659 19864 16635
rect 20911 18734 20987 18768
rect 20911 14676 20987 14710
rect 21415 18734 21491 18768
rect 21415 14676 21491 14710
rect 8073 12135 8107 12311
rect 10141 12135 10175 12311
rect 6073 11172 6107 11548
rect 10131 11172 10165 11548
rect 6185 10086 6219 10562
rect 6723 10086 6757 10562
rect 7121 10086 7155 10562
rect 7659 10086 7693 10562
rect 9051 10104 9085 10580
rect 9589 10104 9623 10580
rect 9983 10104 10017 10580
rect 10521 10104 10555 10580
rect 12033 10677 12067 10853
rect 12191 10677 12225 10853
rect 12349 10677 12383 10853
rect 12507 10677 12541 10853
rect 12665 10677 12699 10853
rect 6185 9044 6219 9520
rect 6723 9044 6757 9520
rect 7121 9044 7155 9520
rect 7659 9044 7693 9520
rect 9051 9019 9085 9495
rect 9589 9019 9623 9495
rect 9983 9019 10017 9495
rect 10521 9019 10555 9495
rect 24843 7911 25619 7945
rect 24843 7653 25619 7687
rect 24843 7205 26519 7239
rect 24843 6947 26519 6981
rect 24843 6689 26519 6723
rect 24843 6431 26519 6465
rect 24843 6173 26519 6207
rect 24843 5915 26519 5949
rect 24843 5657 26519 5691
rect 24843 5399 26519 5433
rect 24843 5141 26519 5175
<< psubdiff >>
rect 2656 42334 2752 42368
rect 2890 42334 3048 42368
rect 3186 42334 3344 42368
rect 3482 42334 3640 42368
rect 3778 42334 3936 42368
rect 4074 42334 4232 42368
rect 4370 42334 4528 42368
rect 4666 42334 4824 42368
rect 4962 42334 5120 42368
rect 5258 42334 5416 42368
rect 5554 42334 5650 42368
rect 2656 42272 2690 42334
rect 2952 42272 2986 42334
rect 2656 36310 2690 36372
rect 3248 42272 3282 42334
rect 2952 36310 2986 36372
rect 3544 42272 3578 42334
rect 3248 36310 3282 36372
rect 3840 42272 3874 42334
rect 3544 36310 3578 36372
rect 4136 42272 4170 42334
rect 3840 36310 3874 36372
rect 4432 42272 4466 42334
rect 4136 36310 4170 36372
rect 4728 42272 4762 42334
rect 4432 36310 4466 36372
rect 5024 42272 5058 42334
rect 4728 36310 4762 36372
rect 5320 42272 5354 42334
rect 5024 36310 5058 36372
rect 5616 42272 5650 42334
rect 5320 36310 5354 36372
rect 5616 36310 5650 36372
rect 2656 36276 2752 36310
rect 2890 36276 3048 36310
rect 3186 36276 3344 36310
rect 3482 36276 3640 36310
rect 3778 36276 3936 36310
rect 4074 36276 4232 36310
rect 4370 36276 4528 36310
rect 4666 36276 4824 36310
rect 4962 36276 5120 36310
rect 5258 36276 5416 36310
rect 5554 36276 5650 36310
rect 2656 36214 2690 36276
rect 2952 36214 2986 36276
rect 2656 30252 2690 30314
rect 3248 36214 3282 36276
rect 2952 30252 2986 30314
rect 3544 36214 3578 36276
rect 3248 30252 3282 30314
rect 3840 36214 3874 36276
rect 3544 30252 3578 30314
rect 4136 36214 4170 36276
rect 3840 30252 3874 30314
rect 4432 36214 4466 36276
rect 4136 30252 4170 30314
rect 4728 36214 4762 36276
rect 4432 30252 4466 30314
rect 5024 36214 5058 36276
rect 4728 30252 4762 30314
rect 5320 36214 5354 36276
rect 5024 30252 5058 30314
rect 5616 36214 5650 36276
rect 5320 30252 5354 30314
rect 5616 30252 5650 30314
rect 2656 30218 2752 30252
rect 2890 30218 3048 30252
rect 3186 30218 3344 30252
rect 3482 30218 3640 30252
rect 3778 30218 3936 30252
rect 4074 30218 4232 30252
rect 4370 30218 4528 30252
rect 4666 30218 4824 30252
rect 4962 30218 5120 30252
rect 5258 30218 5416 30252
rect 5554 30218 5650 30252
rect 7456 28209 7552 28243
rect 10352 28209 10510 28243
rect 13310 28209 13406 28243
rect 7456 28147 7490 28209
rect 10414 28147 10448 28209
rect 7456 27947 7490 28009
rect 13372 28147 13406 28209
rect 10414 27947 10448 28009
rect 13372 27947 13406 28009
rect 7456 27913 7552 27947
rect 10352 27913 10510 27947
rect 13310 27913 13406 27947
rect 7456 27851 7490 27913
rect 10414 27851 10448 27913
rect 7456 27651 7490 27713
rect 13372 27851 13406 27913
rect 10414 27651 10448 27713
rect 13372 27651 13406 27713
rect 7456 27617 7552 27651
rect 10352 27617 10510 27651
rect 13310 27617 13406 27651
rect 7456 27555 7490 27617
rect 10414 27555 10448 27617
rect 7456 27355 7490 27417
rect 13372 27555 13406 27617
rect 10414 27355 10448 27417
rect 13372 27355 13406 27417
rect 7456 27321 7552 27355
rect 10352 27321 10510 27355
rect 13310 27321 13406 27355
rect 7456 27259 7490 27321
rect 10414 27259 10448 27321
rect 7456 27059 7490 27121
rect 13372 27259 13406 27321
rect 10414 27059 10448 27121
rect 13372 27059 13406 27121
rect 7456 27025 7552 27059
rect 10352 27025 10510 27059
rect 13310 27025 13406 27059
rect 7456 26963 7490 27025
rect 10414 26963 10448 27025
rect 7456 26763 7490 26825
rect 13372 26963 13406 27025
rect 13647 28230 14935 28262
rect 13647 28196 13781 28230
rect 13815 28196 13871 28230
rect 13905 28196 13961 28230
rect 13995 28196 14051 28230
rect 14085 28196 14141 28230
rect 14175 28196 14231 28230
rect 14265 28196 14321 28230
rect 14355 28196 14411 28230
rect 14445 28196 14501 28230
rect 14535 28196 14591 28230
rect 14625 28196 14681 28230
rect 14715 28196 14771 28230
rect 14805 28196 14935 28230
rect 13647 28161 14935 28196
rect 13647 28146 13748 28161
rect 13647 28112 13680 28146
rect 13714 28112 13748 28146
rect 13647 28056 13748 28112
rect 14834 28146 14935 28161
rect 14834 28112 14867 28146
rect 14901 28112 14935 28146
rect 13647 28022 13680 28056
rect 13714 28022 13748 28056
rect 13647 27966 13748 28022
rect 13647 27932 13680 27966
rect 13714 27932 13748 27966
rect 13647 27876 13748 27932
rect 13647 27842 13680 27876
rect 13714 27842 13748 27876
rect 13647 27786 13748 27842
rect 13647 27752 13680 27786
rect 13714 27752 13748 27786
rect 13647 27696 13748 27752
rect 13647 27662 13680 27696
rect 13714 27662 13748 27696
rect 13647 27606 13748 27662
rect 13647 27572 13680 27606
rect 13714 27572 13748 27606
rect 13647 27516 13748 27572
rect 13647 27482 13680 27516
rect 13714 27482 13748 27516
rect 13647 27426 13748 27482
rect 13647 27392 13680 27426
rect 13714 27392 13748 27426
rect 13647 27336 13748 27392
rect 13647 27302 13680 27336
rect 13714 27302 13748 27336
rect 13647 27246 13748 27302
rect 13647 27212 13680 27246
rect 13714 27212 13748 27246
rect 13647 27156 13748 27212
rect 13647 27122 13680 27156
rect 13714 27122 13748 27156
rect 14834 28056 14935 28112
rect 14834 28022 14867 28056
rect 14901 28022 14935 28056
rect 14834 27966 14935 28022
rect 14834 27932 14867 27966
rect 14901 27932 14935 27966
rect 14834 27876 14935 27932
rect 14834 27842 14867 27876
rect 14901 27842 14935 27876
rect 14834 27786 14935 27842
rect 14834 27752 14867 27786
rect 14901 27752 14935 27786
rect 14834 27696 14935 27752
rect 14834 27662 14867 27696
rect 14901 27662 14935 27696
rect 14834 27606 14935 27662
rect 14834 27572 14867 27606
rect 14901 27572 14935 27606
rect 14834 27516 14935 27572
rect 14834 27482 14867 27516
rect 14901 27482 14935 27516
rect 14834 27426 14935 27482
rect 14834 27392 14867 27426
rect 14901 27392 14935 27426
rect 14834 27336 14935 27392
rect 14834 27302 14867 27336
rect 14901 27302 14935 27336
rect 14834 27246 14935 27302
rect 14834 27212 14867 27246
rect 14901 27212 14935 27246
rect 14834 27156 14935 27212
rect 13647 27075 13748 27122
rect 14834 27122 14867 27156
rect 14901 27122 14935 27156
rect 14834 27075 14935 27122
rect 13647 27066 14935 27075
rect 13647 27032 13680 27066
rect 13714 27043 14867 27066
rect 13714 27032 13781 27043
rect 13647 27009 13781 27032
rect 13815 27009 13871 27043
rect 13905 27009 13961 27043
rect 13995 27009 14051 27043
rect 14085 27009 14141 27043
rect 14175 27009 14231 27043
rect 14265 27009 14321 27043
rect 14355 27009 14411 27043
rect 14445 27009 14501 27043
rect 14535 27009 14591 27043
rect 14625 27009 14681 27043
rect 14715 27009 14771 27043
rect 14805 27032 14867 27043
rect 14901 27032 14935 27066
rect 14805 27009 14935 27032
rect 13647 26974 14935 27009
rect 14991 28230 16279 28262
rect 14991 28196 15125 28230
rect 15159 28196 15215 28230
rect 15249 28196 15305 28230
rect 15339 28196 15395 28230
rect 15429 28196 15485 28230
rect 15519 28196 15575 28230
rect 15609 28196 15665 28230
rect 15699 28196 15755 28230
rect 15789 28196 15845 28230
rect 15879 28196 15935 28230
rect 15969 28196 16025 28230
rect 16059 28196 16115 28230
rect 16149 28196 16279 28230
rect 14991 28161 16279 28196
rect 14991 28146 15092 28161
rect 14991 28112 15024 28146
rect 15058 28112 15092 28146
rect 14991 28056 15092 28112
rect 16178 28146 16279 28161
rect 16178 28112 16211 28146
rect 16245 28112 16279 28146
rect 14991 28022 15024 28056
rect 15058 28022 15092 28056
rect 14991 27966 15092 28022
rect 14991 27932 15024 27966
rect 15058 27932 15092 27966
rect 14991 27876 15092 27932
rect 14991 27842 15024 27876
rect 15058 27842 15092 27876
rect 14991 27786 15092 27842
rect 14991 27752 15024 27786
rect 15058 27752 15092 27786
rect 14991 27696 15092 27752
rect 14991 27662 15024 27696
rect 15058 27662 15092 27696
rect 14991 27606 15092 27662
rect 14991 27572 15024 27606
rect 15058 27572 15092 27606
rect 14991 27516 15092 27572
rect 14991 27482 15024 27516
rect 15058 27482 15092 27516
rect 14991 27426 15092 27482
rect 14991 27392 15024 27426
rect 15058 27392 15092 27426
rect 14991 27336 15092 27392
rect 14991 27302 15024 27336
rect 15058 27302 15092 27336
rect 14991 27246 15092 27302
rect 14991 27212 15024 27246
rect 15058 27212 15092 27246
rect 14991 27156 15092 27212
rect 14991 27122 15024 27156
rect 15058 27122 15092 27156
rect 16178 28056 16279 28112
rect 16178 28022 16211 28056
rect 16245 28022 16279 28056
rect 16178 27966 16279 28022
rect 16178 27932 16211 27966
rect 16245 27932 16279 27966
rect 16178 27876 16279 27932
rect 16178 27842 16211 27876
rect 16245 27842 16279 27876
rect 16178 27786 16279 27842
rect 16178 27752 16211 27786
rect 16245 27752 16279 27786
rect 16178 27696 16279 27752
rect 16178 27662 16211 27696
rect 16245 27662 16279 27696
rect 16178 27606 16279 27662
rect 16178 27572 16211 27606
rect 16245 27572 16279 27606
rect 16178 27516 16279 27572
rect 16178 27482 16211 27516
rect 16245 27482 16279 27516
rect 16178 27426 16279 27482
rect 16178 27392 16211 27426
rect 16245 27392 16279 27426
rect 16178 27336 16279 27392
rect 16178 27302 16211 27336
rect 16245 27302 16279 27336
rect 16178 27246 16279 27302
rect 16178 27212 16211 27246
rect 16245 27212 16279 27246
rect 16178 27156 16279 27212
rect 14991 27075 15092 27122
rect 16178 27122 16211 27156
rect 16245 27122 16279 27156
rect 16178 27075 16279 27122
rect 14991 27066 16279 27075
rect 14991 27032 15024 27066
rect 15058 27043 16211 27066
rect 15058 27032 15125 27043
rect 14991 27009 15125 27032
rect 15159 27009 15215 27043
rect 15249 27009 15305 27043
rect 15339 27009 15395 27043
rect 15429 27009 15485 27043
rect 15519 27009 15575 27043
rect 15609 27009 15665 27043
rect 15699 27009 15755 27043
rect 15789 27009 15845 27043
rect 15879 27009 15935 27043
rect 15969 27009 16025 27043
rect 16059 27009 16115 27043
rect 16149 27032 16211 27043
rect 16245 27032 16279 27066
rect 16149 27009 16279 27032
rect 14991 26974 16279 27009
rect 16335 28230 17623 28262
rect 16335 28196 16469 28230
rect 16503 28196 16559 28230
rect 16593 28196 16649 28230
rect 16683 28196 16739 28230
rect 16773 28196 16829 28230
rect 16863 28196 16919 28230
rect 16953 28196 17009 28230
rect 17043 28196 17099 28230
rect 17133 28196 17189 28230
rect 17223 28196 17279 28230
rect 17313 28196 17369 28230
rect 17403 28196 17459 28230
rect 17493 28196 17623 28230
rect 16335 28161 17623 28196
rect 16335 28146 16436 28161
rect 16335 28112 16368 28146
rect 16402 28112 16436 28146
rect 16335 28056 16436 28112
rect 17522 28146 17623 28161
rect 17522 28112 17555 28146
rect 17589 28112 17623 28146
rect 16335 28022 16368 28056
rect 16402 28022 16436 28056
rect 16335 27966 16436 28022
rect 16335 27932 16368 27966
rect 16402 27932 16436 27966
rect 16335 27876 16436 27932
rect 16335 27842 16368 27876
rect 16402 27842 16436 27876
rect 16335 27786 16436 27842
rect 16335 27752 16368 27786
rect 16402 27752 16436 27786
rect 16335 27696 16436 27752
rect 16335 27662 16368 27696
rect 16402 27662 16436 27696
rect 16335 27606 16436 27662
rect 16335 27572 16368 27606
rect 16402 27572 16436 27606
rect 16335 27516 16436 27572
rect 16335 27482 16368 27516
rect 16402 27482 16436 27516
rect 16335 27426 16436 27482
rect 16335 27392 16368 27426
rect 16402 27392 16436 27426
rect 16335 27336 16436 27392
rect 16335 27302 16368 27336
rect 16402 27302 16436 27336
rect 16335 27246 16436 27302
rect 16335 27212 16368 27246
rect 16402 27212 16436 27246
rect 16335 27156 16436 27212
rect 16335 27122 16368 27156
rect 16402 27122 16436 27156
rect 17522 28056 17623 28112
rect 17522 28022 17555 28056
rect 17589 28022 17623 28056
rect 17522 27966 17623 28022
rect 17522 27932 17555 27966
rect 17589 27932 17623 27966
rect 17522 27876 17623 27932
rect 17522 27842 17555 27876
rect 17589 27842 17623 27876
rect 17522 27786 17623 27842
rect 17522 27752 17555 27786
rect 17589 27752 17623 27786
rect 17522 27696 17623 27752
rect 17522 27662 17555 27696
rect 17589 27662 17623 27696
rect 17522 27606 17623 27662
rect 17522 27572 17555 27606
rect 17589 27572 17623 27606
rect 17522 27516 17623 27572
rect 17522 27482 17555 27516
rect 17589 27482 17623 27516
rect 17522 27426 17623 27482
rect 17522 27392 17555 27426
rect 17589 27392 17623 27426
rect 17522 27336 17623 27392
rect 17522 27302 17555 27336
rect 17589 27302 17623 27336
rect 17522 27246 17623 27302
rect 17522 27212 17555 27246
rect 17589 27212 17623 27246
rect 17522 27156 17623 27212
rect 16335 27075 16436 27122
rect 17522 27122 17555 27156
rect 17589 27122 17623 27156
rect 17522 27075 17623 27122
rect 16335 27066 17623 27075
rect 16335 27032 16368 27066
rect 16402 27043 17555 27066
rect 16402 27032 16469 27043
rect 16335 27009 16469 27032
rect 16503 27009 16559 27043
rect 16593 27009 16649 27043
rect 16683 27009 16739 27043
rect 16773 27009 16829 27043
rect 16863 27009 16919 27043
rect 16953 27009 17009 27043
rect 17043 27009 17099 27043
rect 17133 27009 17189 27043
rect 17223 27009 17279 27043
rect 17313 27009 17369 27043
rect 17403 27009 17459 27043
rect 17493 27032 17555 27043
rect 17589 27032 17623 27066
rect 17493 27009 17623 27032
rect 16335 26974 17623 27009
rect 10414 26763 10448 26825
rect 13372 26763 13406 26825
rect 7456 26729 7552 26763
rect 10352 26729 10510 26763
rect 13310 26729 13406 26763
rect 7456 26667 7490 26729
rect 10414 26667 10448 26729
rect 7456 26467 7490 26529
rect 13372 26667 13406 26729
rect 10414 26467 10448 26529
rect 13372 26467 13406 26529
rect 7456 26433 7552 26467
rect 10352 26433 10510 26467
rect 13310 26433 13406 26467
rect 7456 26371 7490 26433
rect 10414 26371 10448 26433
rect 7456 26171 7490 26233
rect 13372 26371 13406 26433
rect 10414 26171 10448 26233
rect 13372 26171 13406 26233
rect 7456 26137 7552 26171
rect 10352 26137 10510 26171
rect 13310 26137 13406 26171
rect 7456 26075 7490 26137
rect 10414 26075 10448 26137
rect 7456 25875 7490 25937
rect 13372 26075 13406 26137
rect 10414 25875 10448 25937
rect 13372 25875 13406 25937
rect 7456 25841 7552 25875
rect 10352 25841 10510 25875
rect 13310 25841 13406 25875
rect 7456 25779 7490 25841
rect 10414 25779 10448 25841
rect 7456 25579 7490 25641
rect 13372 25779 13406 25841
rect 10414 25579 10448 25641
rect 13372 25579 13406 25641
rect 13647 26886 14935 26918
rect 13647 26852 13781 26886
rect 13815 26852 13871 26886
rect 13905 26852 13961 26886
rect 13995 26852 14051 26886
rect 14085 26852 14141 26886
rect 14175 26852 14231 26886
rect 14265 26852 14321 26886
rect 14355 26852 14411 26886
rect 14445 26852 14501 26886
rect 14535 26852 14591 26886
rect 14625 26852 14681 26886
rect 14715 26852 14771 26886
rect 14805 26852 14935 26886
rect 13647 26817 14935 26852
rect 13647 26802 13748 26817
rect 13647 26768 13680 26802
rect 13714 26768 13748 26802
rect 13647 26712 13748 26768
rect 14834 26802 14935 26817
rect 14834 26768 14867 26802
rect 14901 26768 14935 26802
rect 13647 26678 13680 26712
rect 13714 26678 13748 26712
rect 13647 26622 13748 26678
rect 13647 26588 13680 26622
rect 13714 26588 13748 26622
rect 13647 26532 13748 26588
rect 13647 26498 13680 26532
rect 13714 26498 13748 26532
rect 13647 26442 13748 26498
rect 13647 26408 13680 26442
rect 13714 26408 13748 26442
rect 13647 26352 13748 26408
rect 13647 26318 13680 26352
rect 13714 26318 13748 26352
rect 13647 26262 13748 26318
rect 13647 26228 13680 26262
rect 13714 26228 13748 26262
rect 13647 26172 13748 26228
rect 13647 26138 13680 26172
rect 13714 26138 13748 26172
rect 13647 26082 13748 26138
rect 13647 26048 13680 26082
rect 13714 26048 13748 26082
rect 13647 25992 13748 26048
rect 13647 25958 13680 25992
rect 13714 25958 13748 25992
rect 13647 25902 13748 25958
rect 13647 25868 13680 25902
rect 13714 25868 13748 25902
rect 13647 25812 13748 25868
rect 13647 25778 13680 25812
rect 13714 25778 13748 25812
rect 14834 26712 14935 26768
rect 14834 26678 14867 26712
rect 14901 26678 14935 26712
rect 14834 26622 14935 26678
rect 14834 26588 14867 26622
rect 14901 26588 14935 26622
rect 14834 26532 14935 26588
rect 14834 26498 14867 26532
rect 14901 26498 14935 26532
rect 14834 26442 14935 26498
rect 14834 26408 14867 26442
rect 14901 26408 14935 26442
rect 14834 26352 14935 26408
rect 14834 26318 14867 26352
rect 14901 26318 14935 26352
rect 14834 26262 14935 26318
rect 14834 26228 14867 26262
rect 14901 26228 14935 26262
rect 14834 26172 14935 26228
rect 14834 26138 14867 26172
rect 14901 26138 14935 26172
rect 14834 26082 14935 26138
rect 14834 26048 14867 26082
rect 14901 26048 14935 26082
rect 14834 25992 14935 26048
rect 14834 25958 14867 25992
rect 14901 25958 14935 25992
rect 14834 25902 14935 25958
rect 14834 25868 14867 25902
rect 14901 25868 14935 25902
rect 14834 25812 14935 25868
rect 13647 25731 13748 25778
rect 14834 25778 14867 25812
rect 14901 25778 14935 25812
rect 14834 25731 14935 25778
rect 13647 25722 14935 25731
rect 13647 25688 13680 25722
rect 13714 25699 14867 25722
rect 13714 25688 13781 25699
rect 13647 25665 13781 25688
rect 13815 25665 13871 25699
rect 13905 25665 13961 25699
rect 13995 25665 14051 25699
rect 14085 25665 14141 25699
rect 14175 25665 14231 25699
rect 14265 25665 14321 25699
rect 14355 25665 14411 25699
rect 14445 25665 14501 25699
rect 14535 25665 14591 25699
rect 14625 25665 14681 25699
rect 14715 25665 14771 25699
rect 14805 25688 14867 25699
rect 14901 25688 14935 25722
rect 14805 25665 14935 25688
rect 13647 25630 14935 25665
rect 14991 26886 16279 26918
rect 14991 26852 15125 26886
rect 15159 26852 15215 26886
rect 15249 26852 15305 26886
rect 15339 26852 15395 26886
rect 15429 26852 15485 26886
rect 15519 26852 15575 26886
rect 15609 26852 15665 26886
rect 15699 26852 15755 26886
rect 15789 26852 15845 26886
rect 15879 26852 15935 26886
rect 15969 26852 16025 26886
rect 16059 26852 16115 26886
rect 16149 26852 16279 26886
rect 14991 26817 16279 26852
rect 14991 26802 15092 26817
rect 14991 26768 15024 26802
rect 15058 26768 15092 26802
rect 14991 26712 15092 26768
rect 16178 26802 16279 26817
rect 16178 26768 16211 26802
rect 16245 26768 16279 26802
rect 14991 26678 15024 26712
rect 15058 26678 15092 26712
rect 14991 26622 15092 26678
rect 14991 26588 15024 26622
rect 15058 26588 15092 26622
rect 14991 26532 15092 26588
rect 14991 26498 15024 26532
rect 15058 26498 15092 26532
rect 14991 26442 15092 26498
rect 14991 26408 15024 26442
rect 15058 26408 15092 26442
rect 14991 26352 15092 26408
rect 14991 26318 15024 26352
rect 15058 26318 15092 26352
rect 14991 26262 15092 26318
rect 14991 26228 15024 26262
rect 15058 26228 15092 26262
rect 14991 26172 15092 26228
rect 14991 26138 15024 26172
rect 15058 26138 15092 26172
rect 14991 26082 15092 26138
rect 14991 26048 15024 26082
rect 15058 26048 15092 26082
rect 14991 25992 15092 26048
rect 14991 25958 15024 25992
rect 15058 25958 15092 25992
rect 14991 25902 15092 25958
rect 14991 25868 15024 25902
rect 15058 25868 15092 25902
rect 14991 25812 15092 25868
rect 14991 25778 15024 25812
rect 15058 25778 15092 25812
rect 16178 26712 16279 26768
rect 16178 26678 16211 26712
rect 16245 26678 16279 26712
rect 16178 26622 16279 26678
rect 16178 26588 16211 26622
rect 16245 26588 16279 26622
rect 16178 26532 16279 26588
rect 16178 26498 16211 26532
rect 16245 26498 16279 26532
rect 16178 26442 16279 26498
rect 16178 26408 16211 26442
rect 16245 26408 16279 26442
rect 16178 26352 16279 26408
rect 16178 26318 16211 26352
rect 16245 26318 16279 26352
rect 16178 26262 16279 26318
rect 16178 26228 16211 26262
rect 16245 26228 16279 26262
rect 16178 26172 16279 26228
rect 16178 26138 16211 26172
rect 16245 26138 16279 26172
rect 16178 26082 16279 26138
rect 16178 26048 16211 26082
rect 16245 26048 16279 26082
rect 16178 25992 16279 26048
rect 16178 25958 16211 25992
rect 16245 25958 16279 25992
rect 16178 25902 16279 25958
rect 16178 25868 16211 25902
rect 16245 25868 16279 25902
rect 16178 25812 16279 25868
rect 14991 25731 15092 25778
rect 16178 25778 16211 25812
rect 16245 25778 16279 25812
rect 16178 25731 16279 25778
rect 14991 25722 16279 25731
rect 14991 25688 15024 25722
rect 15058 25699 16211 25722
rect 15058 25688 15125 25699
rect 14991 25665 15125 25688
rect 15159 25665 15215 25699
rect 15249 25665 15305 25699
rect 15339 25665 15395 25699
rect 15429 25665 15485 25699
rect 15519 25665 15575 25699
rect 15609 25665 15665 25699
rect 15699 25665 15755 25699
rect 15789 25665 15845 25699
rect 15879 25665 15935 25699
rect 15969 25665 16025 25699
rect 16059 25665 16115 25699
rect 16149 25688 16211 25699
rect 16245 25688 16279 25722
rect 16149 25665 16279 25688
rect 14991 25630 16279 25665
rect 16335 26886 17623 26918
rect 16335 26852 16469 26886
rect 16503 26852 16559 26886
rect 16593 26852 16649 26886
rect 16683 26852 16739 26886
rect 16773 26852 16829 26886
rect 16863 26852 16919 26886
rect 16953 26852 17009 26886
rect 17043 26852 17099 26886
rect 17133 26852 17189 26886
rect 17223 26852 17279 26886
rect 17313 26852 17369 26886
rect 17403 26852 17459 26886
rect 17493 26852 17623 26886
rect 16335 26817 17623 26852
rect 16335 26802 16436 26817
rect 16335 26768 16368 26802
rect 16402 26768 16436 26802
rect 16335 26712 16436 26768
rect 17522 26802 17623 26817
rect 17522 26768 17555 26802
rect 17589 26768 17623 26802
rect 16335 26678 16368 26712
rect 16402 26678 16436 26712
rect 16335 26622 16436 26678
rect 16335 26588 16368 26622
rect 16402 26588 16436 26622
rect 16335 26532 16436 26588
rect 16335 26498 16368 26532
rect 16402 26498 16436 26532
rect 16335 26442 16436 26498
rect 16335 26408 16368 26442
rect 16402 26408 16436 26442
rect 16335 26352 16436 26408
rect 16335 26318 16368 26352
rect 16402 26318 16436 26352
rect 16335 26262 16436 26318
rect 16335 26228 16368 26262
rect 16402 26228 16436 26262
rect 16335 26172 16436 26228
rect 16335 26138 16368 26172
rect 16402 26138 16436 26172
rect 16335 26082 16436 26138
rect 16335 26048 16368 26082
rect 16402 26048 16436 26082
rect 16335 25992 16436 26048
rect 16335 25958 16368 25992
rect 16402 25958 16436 25992
rect 16335 25902 16436 25958
rect 16335 25868 16368 25902
rect 16402 25868 16436 25902
rect 16335 25812 16436 25868
rect 16335 25778 16368 25812
rect 16402 25778 16436 25812
rect 17522 26712 17623 26768
rect 17522 26678 17555 26712
rect 17589 26678 17623 26712
rect 17522 26622 17623 26678
rect 17522 26588 17555 26622
rect 17589 26588 17623 26622
rect 17522 26532 17623 26588
rect 17522 26498 17555 26532
rect 17589 26498 17623 26532
rect 17522 26442 17623 26498
rect 17522 26408 17555 26442
rect 17589 26408 17623 26442
rect 17522 26352 17623 26408
rect 17522 26318 17555 26352
rect 17589 26318 17623 26352
rect 17522 26262 17623 26318
rect 17522 26228 17555 26262
rect 17589 26228 17623 26262
rect 17522 26172 17623 26228
rect 17522 26138 17555 26172
rect 17589 26138 17623 26172
rect 17522 26082 17623 26138
rect 17522 26048 17555 26082
rect 17589 26048 17623 26082
rect 17522 25992 17623 26048
rect 17522 25958 17555 25992
rect 17589 25958 17623 25992
rect 17522 25902 17623 25958
rect 17522 25868 17555 25902
rect 17589 25868 17623 25902
rect 17522 25812 17623 25868
rect 16335 25731 16436 25778
rect 17522 25778 17555 25812
rect 17589 25778 17623 25812
rect 17522 25731 17623 25778
rect 16335 25722 17623 25731
rect 16335 25688 16368 25722
rect 16402 25699 17555 25722
rect 16402 25688 16469 25699
rect 16335 25665 16469 25688
rect 16503 25665 16559 25699
rect 16593 25665 16649 25699
rect 16683 25665 16739 25699
rect 16773 25665 16829 25699
rect 16863 25665 16919 25699
rect 16953 25665 17009 25699
rect 17043 25665 17099 25699
rect 17133 25665 17189 25699
rect 17223 25665 17279 25699
rect 17313 25665 17369 25699
rect 17403 25665 17459 25699
rect 17493 25688 17555 25699
rect 17589 25688 17623 25722
rect 17493 25665 17623 25688
rect 16335 25630 17623 25665
rect 7456 25545 7552 25579
rect 10352 25545 10510 25579
rect 13310 25545 13406 25579
rect 7456 25483 7490 25545
rect 10414 25483 10448 25545
rect 7456 25283 7490 25345
rect 13372 25483 13406 25545
rect 10414 25283 10448 25345
rect 13372 25283 13406 25345
rect 7456 25249 7552 25283
rect 10352 25249 10510 25283
rect 13310 25249 13406 25283
rect 7456 25187 7490 25249
rect 10414 25187 10448 25249
rect 7456 24987 7490 25049
rect 13372 25187 13406 25249
rect 10414 24987 10448 25049
rect 13372 24987 13406 25049
rect 7456 24953 7552 24987
rect 10352 24953 10510 24987
rect 13310 24953 13406 24987
rect 7456 24891 7490 24953
rect 10414 24891 10448 24953
rect 7456 24691 7490 24753
rect 13372 24891 13406 24953
rect 10414 24691 10448 24753
rect 13372 24691 13406 24753
rect 7456 24657 7552 24691
rect 10352 24657 10510 24691
rect 13310 24657 13406 24691
rect 13647 25542 14935 25574
rect 13647 25508 13781 25542
rect 13815 25508 13871 25542
rect 13905 25508 13961 25542
rect 13995 25508 14051 25542
rect 14085 25508 14141 25542
rect 14175 25508 14231 25542
rect 14265 25508 14321 25542
rect 14355 25508 14411 25542
rect 14445 25508 14501 25542
rect 14535 25508 14591 25542
rect 14625 25508 14681 25542
rect 14715 25508 14771 25542
rect 14805 25508 14935 25542
rect 13647 25473 14935 25508
rect 13647 25458 13748 25473
rect 13647 25424 13680 25458
rect 13714 25424 13748 25458
rect 13647 25368 13748 25424
rect 14834 25458 14935 25473
rect 14834 25424 14867 25458
rect 14901 25424 14935 25458
rect 13647 25334 13680 25368
rect 13714 25334 13748 25368
rect 13647 25278 13748 25334
rect 13647 25244 13680 25278
rect 13714 25244 13748 25278
rect 13647 25188 13748 25244
rect 13647 25154 13680 25188
rect 13714 25154 13748 25188
rect 13647 25098 13748 25154
rect 13647 25064 13680 25098
rect 13714 25064 13748 25098
rect 13647 25008 13748 25064
rect 13647 24974 13680 25008
rect 13714 24974 13748 25008
rect 13647 24918 13748 24974
rect 13647 24884 13680 24918
rect 13714 24884 13748 24918
rect 13647 24828 13748 24884
rect 13647 24794 13680 24828
rect 13714 24794 13748 24828
rect 13647 24738 13748 24794
rect 13647 24704 13680 24738
rect 13714 24704 13748 24738
rect 13647 24648 13748 24704
rect 13647 24614 13680 24648
rect 13714 24614 13748 24648
rect 13647 24558 13748 24614
rect 13647 24524 13680 24558
rect 13714 24524 13748 24558
rect 13647 24468 13748 24524
rect 13647 24434 13680 24468
rect 13714 24434 13748 24468
rect 14834 25368 14935 25424
rect 14834 25334 14867 25368
rect 14901 25334 14935 25368
rect 14834 25278 14935 25334
rect 14834 25244 14867 25278
rect 14901 25244 14935 25278
rect 14834 25188 14935 25244
rect 14834 25154 14867 25188
rect 14901 25154 14935 25188
rect 14834 25098 14935 25154
rect 14834 25064 14867 25098
rect 14901 25064 14935 25098
rect 14834 25008 14935 25064
rect 14834 24974 14867 25008
rect 14901 24974 14935 25008
rect 14834 24918 14935 24974
rect 14834 24884 14867 24918
rect 14901 24884 14935 24918
rect 14834 24828 14935 24884
rect 14834 24794 14867 24828
rect 14901 24794 14935 24828
rect 14834 24738 14935 24794
rect 14834 24704 14867 24738
rect 14901 24704 14935 24738
rect 14834 24648 14935 24704
rect 14834 24614 14867 24648
rect 14901 24614 14935 24648
rect 14834 24558 14935 24614
rect 14834 24524 14867 24558
rect 14901 24524 14935 24558
rect 14834 24468 14935 24524
rect 13647 24387 13748 24434
rect 14834 24434 14867 24468
rect 14901 24434 14935 24468
rect 14834 24387 14935 24434
rect 13647 24378 14935 24387
rect 13647 24344 13680 24378
rect 13714 24355 14867 24378
rect 13714 24344 13781 24355
rect 13647 24321 13781 24344
rect 13815 24321 13871 24355
rect 13905 24321 13961 24355
rect 13995 24321 14051 24355
rect 14085 24321 14141 24355
rect 14175 24321 14231 24355
rect 14265 24321 14321 24355
rect 14355 24321 14411 24355
rect 14445 24321 14501 24355
rect 14535 24321 14591 24355
rect 14625 24321 14681 24355
rect 14715 24321 14771 24355
rect 14805 24344 14867 24355
rect 14901 24344 14935 24378
rect 14805 24321 14935 24344
rect 13647 24286 14935 24321
rect 14991 25542 16279 25574
rect 14991 25508 15125 25542
rect 15159 25508 15215 25542
rect 15249 25508 15305 25542
rect 15339 25508 15395 25542
rect 15429 25508 15485 25542
rect 15519 25508 15575 25542
rect 15609 25508 15665 25542
rect 15699 25508 15755 25542
rect 15789 25508 15845 25542
rect 15879 25508 15935 25542
rect 15969 25508 16025 25542
rect 16059 25508 16115 25542
rect 16149 25508 16279 25542
rect 14991 25473 16279 25508
rect 14991 25458 15092 25473
rect 14991 25424 15024 25458
rect 15058 25424 15092 25458
rect 14991 25368 15092 25424
rect 16178 25458 16279 25473
rect 16178 25424 16211 25458
rect 16245 25424 16279 25458
rect 14991 25334 15024 25368
rect 15058 25334 15092 25368
rect 14991 25278 15092 25334
rect 14991 25244 15024 25278
rect 15058 25244 15092 25278
rect 14991 25188 15092 25244
rect 14991 25154 15024 25188
rect 15058 25154 15092 25188
rect 14991 25098 15092 25154
rect 14991 25064 15024 25098
rect 15058 25064 15092 25098
rect 14991 25008 15092 25064
rect 14991 24974 15024 25008
rect 15058 24974 15092 25008
rect 14991 24918 15092 24974
rect 14991 24884 15024 24918
rect 15058 24884 15092 24918
rect 14991 24828 15092 24884
rect 14991 24794 15024 24828
rect 15058 24794 15092 24828
rect 14991 24738 15092 24794
rect 14991 24704 15024 24738
rect 15058 24704 15092 24738
rect 14991 24648 15092 24704
rect 14991 24614 15024 24648
rect 15058 24614 15092 24648
rect 14991 24558 15092 24614
rect 14991 24524 15024 24558
rect 15058 24524 15092 24558
rect 14991 24468 15092 24524
rect 14991 24434 15024 24468
rect 15058 24434 15092 24468
rect 16178 25368 16279 25424
rect 16178 25334 16211 25368
rect 16245 25334 16279 25368
rect 16178 25278 16279 25334
rect 16178 25244 16211 25278
rect 16245 25244 16279 25278
rect 16178 25188 16279 25244
rect 16178 25154 16211 25188
rect 16245 25154 16279 25188
rect 16178 25098 16279 25154
rect 16178 25064 16211 25098
rect 16245 25064 16279 25098
rect 16178 25008 16279 25064
rect 16178 24974 16211 25008
rect 16245 24974 16279 25008
rect 16178 24918 16279 24974
rect 16178 24884 16211 24918
rect 16245 24884 16279 24918
rect 16178 24828 16279 24884
rect 16178 24794 16211 24828
rect 16245 24794 16279 24828
rect 16178 24738 16279 24794
rect 16178 24704 16211 24738
rect 16245 24704 16279 24738
rect 16178 24648 16279 24704
rect 16178 24614 16211 24648
rect 16245 24614 16279 24648
rect 16178 24558 16279 24614
rect 16178 24524 16211 24558
rect 16245 24524 16279 24558
rect 16178 24468 16279 24524
rect 14991 24387 15092 24434
rect 16178 24434 16211 24468
rect 16245 24434 16279 24468
rect 16178 24387 16279 24434
rect 14991 24378 16279 24387
rect 14991 24344 15024 24378
rect 15058 24355 16211 24378
rect 15058 24344 15125 24355
rect 14991 24321 15125 24344
rect 15159 24321 15215 24355
rect 15249 24321 15305 24355
rect 15339 24321 15395 24355
rect 15429 24321 15485 24355
rect 15519 24321 15575 24355
rect 15609 24321 15665 24355
rect 15699 24321 15755 24355
rect 15789 24321 15845 24355
rect 15879 24321 15935 24355
rect 15969 24321 16025 24355
rect 16059 24321 16115 24355
rect 16149 24344 16211 24355
rect 16245 24344 16279 24378
rect 16149 24321 16279 24344
rect 14991 24286 16279 24321
rect 16335 25542 17623 25574
rect 16335 25508 16469 25542
rect 16503 25508 16559 25542
rect 16593 25508 16649 25542
rect 16683 25508 16739 25542
rect 16773 25508 16829 25542
rect 16863 25508 16919 25542
rect 16953 25508 17009 25542
rect 17043 25508 17099 25542
rect 17133 25508 17189 25542
rect 17223 25508 17279 25542
rect 17313 25508 17369 25542
rect 17403 25508 17459 25542
rect 17493 25508 17623 25542
rect 16335 25473 17623 25508
rect 16335 25458 16436 25473
rect 16335 25424 16368 25458
rect 16402 25424 16436 25458
rect 16335 25368 16436 25424
rect 17522 25458 17623 25473
rect 17522 25424 17555 25458
rect 17589 25424 17623 25458
rect 16335 25334 16368 25368
rect 16402 25334 16436 25368
rect 16335 25278 16436 25334
rect 16335 25244 16368 25278
rect 16402 25244 16436 25278
rect 16335 25188 16436 25244
rect 16335 25154 16368 25188
rect 16402 25154 16436 25188
rect 16335 25098 16436 25154
rect 16335 25064 16368 25098
rect 16402 25064 16436 25098
rect 16335 25008 16436 25064
rect 16335 24974 16368 25008
rect 16402 24974 16436 25008
rect 16335 24918 16436 24974
rect 16335 24884 16368 24918
rect 16402 24884 16436 24918
rect 16335 24828 16436 24884
rect 16335 24794 16368 24828
rect 16402 24794 16436 24828
rect 16335 24738 16436 24794
rect 16335 24704 16368 24738
rect 16402 24704 16436 24738
rect 16335 24648 16436 24704
rect 16335 24614 16368 24648
rect 16402 24614 16436 24648
rect 16335 24558 16436 24614
rect 16335 24524 16368 24558
rect 16402 24524 16436 24558
rect 16335 24468 16436 24524
rect 16335 24434 16368 24468
rect 16402 24434 16436 24468
rect 17522 25368 17623 25424
rect 17522 25334 17555 25368
rect 17589 25334 17623 25368
rect 17522 25278 17623 25334
rect 17522 25244 17555 25278
rect 17589 25244 17623 25278
rect 17522 25188 17623 25244
rect 17522 25154 17555 25188
rect 17589 25154 17623 25188
rect 17522 25098 17623 25154
rect 17522 25064 17555 25098
rect 17589 25064 17623 25098
rect 17522 25008 17623 25064
rect 17522 24974 17555 25008
rect 17589 24974 17623 25008
rect 17522 24918 17623 24974
rect 17522 24884 17555 24918
rect 17589 24884 17623 24918
rect 17522 24828 17623 24884
rect 17522 24794 17555 24828
rect 17589 24794 17623 24828
rect 17522 24738 17623 24794
rect 17522 24704 17555 24738
rect 17589 24704 17623 24738
rect 17522 24648 17623 24704
rect 17522 24614 17555 24648
rect 17589 24614 17623 24648
rect 17522 24558 17623 24614
rect 17522 24524 17555 24558
rect 17589 24524 17623 24558
rect 17522 24468 17623 24524
rect 16335 24387 16436 24434
rect 17522 24434 17555 24468
rect 17589 24434 17623 24468
rect 17522 24387 17623 24434
rect 16335 24378 17623 24387
rect 16335 24344 16368 24378
rect 16402 24355 17555 24378
rect 16402 24344 16469 24355
rect 16335 24321 16469 24344
rect 16503 24321 16559 24355
rect 16593 24321 16649 24355
rect 16683 24321 16739 24355
rect 16773 24321 16829 24355
rect 16863 24321 16919 24355
rect 16953 24321 17009 24355
rect 17043 24321 17099 24355
rect 17133 24321 17189 24355
rect 17223 24321 17279 24355
rect 17313 24321 17369 24355
rect 17403 24321 17459 24355
rect 17493 24344 17555 24355
rect 17589 24344 17623 24378
rect 17493 24321 17623 24344
rect 16335 24286 17623 24321
rect 13967 10793 14063 10827
rect 14201 10793 14359 10827
rect 14497 10793 14655 10827
rect 14793 10793 14951 10827
rect 15089 10793 15247 10827
rect 15385 10793 15543 10827
rect 15681 10793 15839 10827
rect 15977 10793 16135 10827
rect 16273 10793 16369 10827
rect 13967 10731 14001 10793
rect 14263 10731 14297 10793
rect 13967 6669 14001 6731
rect 14559 10731 14593 10793
rect 14263 6669 14297 6731
rect 14855 10731 14889 10793
rect 14559 6669 14593 6731
rect 15151 10731 15185 10793
rect 14855 6669 14889 6731
rect 15447 10731 15481 10793
rect 15151 6669 15185 6731
rect 15743 10731 15777 10793
rect 15447 6669 15481 6731
rect 16039 10731 16073 10793
rect 15743 6669 15777 6731
rect 16335 10731 16369 10793
rect 16039 6669 16073 6731
rect 16335 6669 16369 6731
rect 13967 6635 14063 6669
rect 14201 6635 14359 6669
rect 14497 6635 14655 6669
rect 14793 6635 14951 6669
rect 15089 6635 15247 6669
rect 15385 6635 15543 6669
rect 15681 6635 15839 6669
rect 15977 6635 16135 6669
rect 16273 6635 16369 6669
rect 13967 6573 14001 6635
rect 14263 6573 14297 6635
rect 13967 2511 14001 2573
rect 14559 6573 14593 6635
rect 14263 2511 14297 2573
rect 14855 6573 14889 6635
rect 14559 2511 14593 2573
rect 15151 6573 15185 6635
rect 14855 2511 14889 2573
rect 15447 6573 15481 6635
rect 15151 2511 15185 2573
rect 15743 6573 15777 6635
rect 15447 2511 15481 2573
rect 16039 6573 16073 6635
rect 15743 2511 15777 2573
rect 16335 6573 16369 6635
rect 16039 2511 16073 2573
rect 18584 6335 18680 6369
rect 18818 6335 18976 6369
rect 19114 6335 19272 6369
rect 19410 6335 19568 6369
rect 19706 6335 19802 6369
rect 18584 6273 18618 6335
rect 16335 2511 16369 2573
rect 13967 2477 14063 2511
rect 14201 2477 14359 2511
rect 14497 2477 14655 2511
rect 14793 2477 14951 2511
rect 15089 2477 15247 2511
rect 15385 2477 15543 2511
rect 15681 2477 15839 2511
rect 15977 2477 16135 2511
rect 16273 2477 16369 2511
rect 18880 6273 18914 6335
rect 18584 2511 18618 2573
rect 19176 6273 19210 6335
rect 18880 2511 18914 2573
rect 19472 6273 19506 6335
rect 19176 2511 19210 2573
rect 19768 6273 19802 6335
rect 19472 2511 19506 2573
rect 19768 2511 19802 2573
rect 18584 2477 18680 2511
rect 18818 2477 18976 2511
rect 19114 2477 19272 2511
rect 19410 2477 19568 2511
rect 19706 2477 19802 2511
<< nsubdiff >>
rect 13810 28080 14772 28099
rect 13810 28046 13921 28080
rect 13955 28046 14011 28080
rect 14045 28046 14101 28080
rect 14135 28046 14191 28080
rect 14225 28046 14281 28080
rect 14315 28046 14371 28080
rect 14405 28046 14461 28080
rect 14495 28046 14551 28080
rect 14585 28046 14641 28080
rect 14675 28046 14772 28080
rect 13810 28027 14772 28046
rect 13810 27986 13882 28027
rect 13810 27952 13829 27986
rect 13863 27952 13882 27986
rect 14700 27967 14772 28027
rect 13810 27896 13882 27952
rect 13810 27862 13829 27896
rect 13863 27862 13882 27896
rect 13810 27806 13882 27862
rect 13810 27772 13829 27806
rect 13863 27772 13882 27806
rect 13810 27716 13882 27772
rect 13810 27682 13829 27716
rect 13863 27682 13882 27716
rect 13810 27626 13882 27682
rect 13810 27592 13829 27626
rect 13863 27592 13882 27626
rect 13810 27536 13882 27592
rect 13810 27502 13829 27536
rect 13863 27502 13882 27536
rect 13810 27446 13882 27502
rect 13810 27412 13829 27446
rect 13863 27412 13882 27446
rect 13810 27356 13882 27412
rect 13810 27322 13829 27356
rect 13863 27322 13882 27356
rect 13810 27266 13882 27322
rect 14700 27933 14719 27967
rect 14753 27933 14772 27967
rect 14700 27877 14772 27933
rect 14700 27843 14719 27877
rect 14753 27843 14772 27877
rect 14700 27787 14772 27843
rect 14700 27753 14719 27787
rect 14753 27753 14772 27787
rect 14700 27697 14772 27753
rect 14700 27663 14719 27697
rect 14753 27663 14772 27697
rect 14700 27607 14772 27663
rect 14700 27573 14719 27607
rect 14753 27573 14772 27607
rect 14700 27517 14772 27573
rect 14700 27483 14719 27517
rect 14753 27483 14772 27517
rect 14700 27427 14772 27483
rect 14700 27393 14719 27427
rect 14753 27393 14772 27427
rect 14700 27337 14772 27393
rect 14700 27303 14719 27337
rect 14753 27303 14772 27337
rect 13810 27232 13829 27266
rect 13863 27232 13882 27266
rect 13810 27209 13882 27232
rect 14700 27247 14772 27303
rect 14700 27213 14719 27247
rect 14753 27213 14772 27247
rect 14700 27209 14772 27213
rect 13810 27190 14772 27209
rect 13810 27156 13887 27190
rect 13921 27156 13977 27190
rect 14011 27156 14067 27190
rect 14101 27156 14157 27190
rect 14191 27156 14247 27190
rect 14281 27156 14337 27190
rect 14371 27156 14427 27190
rect 14461 27156 14517 27190
rect 14551 27156 14607 27190
rect 14641 27156 14772 27190
rect 13810 27137 14772 27156
rect 15154 28080 16116 28099
rect 15154 28046 15265 28080
rect 15299 28046 15355 28080
rect 15389 28046 15445 28080
rect 15479 28046 15535 28080
rect 15569 28046 15625 28080
rect 15659 28046 15715 28080
rect 15749 28046 15805 28080
rect 15839 28046 15895 28080
rect 15929 28046 15985 28080
rect 16019 28046 16116 28080
rect 15154 28027 16116 28046
rect 15154 27986 15226 28027
rect 15154 27952 15173 27986
rect 15207 27952 15226 27986
rect 16044 27967 16116 28027
rect 15154 27896 15226 27952
rect 15154 27862 15173 27896
rect 15207 27862 15226 27896
rect 15154 27806 15226 27862
rect 15154 27772 15173 27806
rect 15207 27772 15226 27806
rect 15154 27716 15226 27772
rect 15154 27682 15173 27716
rect 15207 27682 15226 27716
rect 15154 27626 15226 27682
rect 15154 27592 15173 27626
rect 15207 27592 15226 27626
rect 15154 27536 15226 27592
rect 15154 27502 15173 27536
rect 15207 27502 15226 27536
rect 15154 27446 15226 27502
rect 15154 27412 15173 27446
rect 15207 27412 15226 27446
rect 15154 27356 15226 27412
rect 15154 27322 15173 27356
rect 15207 27322 15226 27356
rect 15154 27266 15226 27322
rect 16044 27933 16063 27967
rect 16097 27933 16116 27967
rect 16044 27877 16116 27933
rect 16044 27843 16063 27877
rect 16097 27843 16116 27877
rect 16044 27787 16116 27843
rect 16044 27753 16063 27787
rect 16097 27753 16116 27787
rect 16044 27697 16116 27753
rect 16044 27663 16063 27697
rect 16097 27663 16116 27697
rect 16044 27607 16116 27663
rect 16044 27573 16063 27607
rect 16097 27573 16116 27607
rect 16044 27517 16116 27573
rect 16044 27483 16063 27517
rect 16097 27483 16116 27517
rect 16044 27427 16116 27483
rect 16044 27393 16063 27427
rect 16097 27393 16116 27427
rect 16044 27337 16116 27393
rect 16044 27303 16063 27337
rect 16097 27303 16116 27337
rect 15154 27232 15173 27266
rect 15207 27232 15226 27266
rect 15154 27209 15226 27232
rect 16044 27247 16116 27303
rect 16044 27213 16063 27247
rect 16097 27213 16116 27247
rect 16044 27209 16116 27213
rect 15154 27190 16116 27209
rect 15154 27156 15231 27190
rect 15265 27156 15321 27190
rect 15355 27156 15411 27190
rect 15445 27156 15501 27190
rect 15535 27156 15591 27190
rect 15625 27156 15681 27190
rect 15715 27156 15771 27190
rect 15805 27156 15861 27190
rect 15895 27156 15951 27190
rect 15985 27156 16116 27190
rect 15154 27137 16116 27156
rect 16498 28080 17460 28099
rect 16498 28046 16609 28080
rect 16643 28046 16699 28080
rect 16733 28046 16789 28080
rect 16823 28046 16879 28080
rect 16913 28046 16969 28080
rect 17003 28046 17059 28080
rect 17093 28046 17149 28080
rect 17183 28046 17239 28080
rect 17273 28046 17329 28080
rect 17363 28046 17460 28080
rect 16498 28027 17460 28046
rect 16498 27986 16570 28027
rect 16498 27952 16517 27986
rect 16551 27952 16570 27986
rect 17388 27967 17460 28027
rect 16498 27896 16570 27952
rect 16498 27862 16517 27896
rect 16551 27862 16570 27896
rect 16498 27806 16570 27862
rect 16498 27772 16517 27806
rect 16551 27772 16570 27806
rect 16498 27716 16570 27772
rect 16498 27682 16517 27716
rect 16551 27682 16570 27716
rect 16498 27626 16570 27682
rect 16498 27592 16517 27626
rect 16551 27592 16570 27626
rect 16498 27536 16570 27592
rect 16498 27502 16517 27536
rect 16551 27502 16570 27536
rect 16498 27446 16570 27502
rect 16498 27412 16517 27446
rect 16551 27412 16570 27446
rect 16498 27356 16570 27412
rect 16498 27322 16517 27356
rect 16551 27322 16570 27356
rect 16498 27266 16570 27322
rect 17388 27933 17407 27967
rect 17441 27933 17460 27967
rect 17388 27877 17460 27933
rect 17388 27843 17407 27877
rect 17441 27843 17460 27877
rect 17388 27787 17460 27843
rect 17388 27753 17407 27787
rect 17441 27753 17460 27787
rect 17388 27697 17460 27753
rect 17388 27663 17407 27697
rect 17441 27663 17460 27697
rect 17388 27607 17460 27663
rect 17388 27573 17407 27607
rect 17441 27573 17460 27607
rect 17388 27517 17460 27573
rect 17388 27483 17407 27517
rect 17441 27483 17460 27517
rect 17388 27427 17460 27483
rect 17388 27393 17407 27427
rect 17441 27393 17460 27427
rect 17388 27337 17460 27393
rect 17388 27303 17407 27337
rect 17441 27303 17460 27337
rect 16498 27232 16517 27266
rect 16551 27232 16570 27266
rect 16498 27209 16570 27232
rect 17388 27247 17460 27303
rect 17388 27213 17407 27247
rect 17441 27213 17460 27247
rect 17388 27209 17460 27213
rect 16498 27190 17460 27209
rect 16498 27156 16575 27190
rect 16609 27156 16665 27190
rect 16699 27156 16755 27190
rect 16789 27156 16845 27190
rect 16879 27156 16935 27190
rect 16969 27156 17025 27190
rect 17059 27156 17115 27190
rect 17149 27156 17205 27190
rect 17239 27156 17295 27190
rect 17329 27156 17460 27190
rect 16498 27137 17460 27156
rect 13810 26736 14772 26755
rect 13810 26702 13921 26736
rect 13955 26702 14011 26736
rect 14045 26702 14101 26736
rect 14135 26702 14191 26736
rect 14225 26702 14281 26736
rect 14315 26702 14371 26736
rect 14405 26702 14461 26736
rect 14495 26702 14551 26736
rect 14585 26702 14641 26736
rect 14675 26702 14772 26736
rect 13810 26683 14772 26702
rect 13810 26642 13882 26683
rect 13810 26608 13829 26642
rect 13863 26608 13882 26642
rect 14700 26623 14772 26683
rect 13810 26552 13882 26608
rect 13810 26518 13829 26552
rect 13863 26518 13882 26552
rect 13810 26462 13882 26518
rect 13810 26428 13829 26462
rect 13863 26428 13882 26462
rect 13810 26372 13882 26428
rect 13810 26338 13829 26372
rect 13863 26338 13882 26372
rect 13810 26282 13882 26338
rect 13810 26248 13829 26282
rect 13863 26248 13882 26282
rect 13810 26192 13882 26248
rect 13810 26158 13829 26192
rect 13863 26158 13882 26192
rect 13810 26102 13882 26158
rect 13810 26068 13829 26102
rect 13863 26068 13882 26102
rect 13810 26012 13882 26068
rect 13810 25978 13829 26012
rect 13863 25978 13882 26012
rect 13810 25922 13882 25978
rect 14700 26589 14719 26623
rect 14753 26589 14772 26623
rect 14700 26533 14772 26589
rect 14700 26499 14719 26533
rect 14753 26499 14772 26533
rect 14700 26443 14772 26499
rect 14700 26409 14719 26443
rect 14753 26409 14772 26443
rect 14700 26353 14772 26409
rect 14700 26319 14719 26353
rect 14753 26319 14772 26353
rect 14700 26263 14772 26319
rect 14700 26229 14719 26263
rect 14753 26229 14772 26263
rect 14700 26173 14772 26229
rect 14700 26139 14719 26173
rect 14753 26139 14772 26173
rect 14700 26083 14772 26139
rect 14700 26049 14719 26083
rect 14753 26049 14772 26083
rect 14700 25993 14772 26049
rect 14700 25959 14719 25993
rect 14753 25959 14772 25993
rect 13810 25888 13829 25922
rect 13863 25888 13882 25922
rect 13810 25865 13882 25888
rect 14700 25903 14772 25959
rect 14700 25869 14719 25903
rect 14753 25869 14772 25903
rect 14700 25865 14772 25869
rect 13810 25846 14772 25865
rect 13810 25812 13887 25846
rect 13921 25812 13977 25846
rect 14011 25812 14067 25846
rect 14101 25812 14157 25846
rect 14191 25812 14247 25846
rect 14281 25812 14337 25846
rect 14371 25812 14427 25846
rect 14461 25812 14517 25846
rect 14551 25812 14607 25846
rect 14641 25812 14772 25846
rect 13810 25793 14772 25812
rect 15154 26736 16116 26755
rect 15154 26702 15265 26736
rect 15299 26702 15355 26736
rect 15389 26702 15445 26736
rect 15479 26702 15535 26736
rect 15569 26702 15625 26736
rect 15659 26702 15715 26736
rect 15749 26702 15805 26736
rect 15839 26702 15895 26736
rect 15929 26702 15985 26736
rect 16019 26702 16116 26736
rect 15154 26683 16116 26702
rect 15154 26642 15226 26683
rect 15154 26608 15173 26642
rect 15207 26608 15226 26642
rect 16044 26623 16116 26683
rect 15154 26552 15226 26608
rect 15154 26518 15173 26552
rect 15207 26518 15226 26552
rect 15154 26462 15226 26518
rect 15154 26428 15173 26462
rect 15207 26428 15226 26462
rect 15154 26372 15226 26428
rect 15154 26338 15173 26372
rect 15207 26338 15226 26372
rect 15154 26282 15226 26338
rect 15154 26248 15173 26282
rect 15207 26248 15226 26282
rect 15154 26192 15226 26248
rect 15154 26158 15173 26192
rect 15207 26158 15226 26192
rect 15154 26102 15226 26158
rect 15154 26068 15173 26102
rect 15207 26068 15226 26102
rect 15154 26012 15226 26068
rect 15154 25978 15173 26012
rect 15207 25978 15226 26012
rect 15154 25922 15226 25978
rect 16044 26589 16063 26623
rect 16097 26589 16116 26623
rect 16044 26533 16116 26589
rect 16044 26499 16063 26533
rect 16097 26499 16116 26533
rect 16044 26443 16116 26499
rect 16044 26409 16063 26443
rect 16097 26409 16116 26443
rect 16044 26353 16116 26409
rect 16044 26319 16063 26353
rect 16097 26319 16116 26353
rect 16044 26263 16116 26319
rect 16044 26229 16063 26263
rect 16097 26229 16116 26263
rect 16044 26173 16116 26229
rect 16044 26139 16063 26173
rect 16097 26139 16116 26173
rect 16044 26083 16116 26139
rect 16044 26049 16063 26083
rect 16097 26049 16116 26083
rect 16044 25993 16116 26049
rect 16044 25959 16063 25993
rect 16097 25959 16116 25993
rect 15154 25888 15173 25922
rect 15207 25888 15226 25922
rect 15154 25865 15226 25888
rect 16044 25903 16116 25959
rect 16044 25869 16063 25903
rect 16097 25869 16116 25903
rect 16044 25865 16116 25869
rect 15154 25846 16116 25865
rect 15154 25812 15231 25846
rect 15265 25812 15321 25846
rect 15355 25812 15411 25846
rect 15445 25812 15501 25846
rect 15535 25812 15591 25846
rect 15625 25812 15681 25846
rect 15715 25812 15771 25846
rect 15805 25812 15861 25846
rect 15895 25812 15951 25846
rect 15985 25812 16116 25846
rect 15154 25793 16116 25812
rect 16498 26736 17460 26755
rect 16498 26702 16609 26736
rect 16643 26702 16699 26736
rect 16733 26702 16789 26736
rect 16823 26702 16879 26736
rect 16913 26702 16969 26736
rect 17003 26702 17059 26736
rect 17093 26702 17149 26736
rect 17183 26702 17239 26736
rect 17273 26702 17329 26736
rect 17363 26702 17460 26736
rect 16498 26683 17460 26702
rect 16498 26642 16570 26683
rect 16498 26608 16517 26642
rect 16551 26608 16570 26642
rect 17388 26623 17460 26683
rect 16498 26552 16570 26608
rect 16498 26518 16517 26552
rect 16551 26518 16570 26552
rect 16498 26462 16570 26518
rect 16498 26428 16517 26462
rect 16551 26428 16570 26462
rect 16498 26372 16570 26428
rect 16498 26338 16517 26372
rect 16551 26338 16570 26372
rect 16498 26282 16570 26338
rect 16498 26248 16517 26282
rect 16551 26248 16570 26282
rect 16498 26192 16570 26248
rect 16498 26158 16517 26192
rect 16551 26158 16570 26192
rect 16498 26102 16570 26158
rect 16498 26068 16517 26102
rect 16551 26068 16570 26102
rect 16498 26012 16570 26068
rect 16498 25978 16517 26012
rect 16551 25978 16570 26012
rect 16498 25922 16570 25978
rect 17388 26589 17407 26623
rect 17441 26589 17460 26623
rect 17388 26533 17460 26589
rect 17388 26499 17407 26533
rect 17441 26499 17460 26533
rect 17388 26443 17460 26499
rect 17388 26409 17407 26443
rect 17441 26409 17460 26443
rect 17388 26353 17460 26409
rect 17388 26319 17407 26353
rect 17441 26319 17460 26353
rect 17388 26263 17460 26319
rect 17388 26229 17407 26263
rect 17441 26229 17460 26263
rect 17388 26173 17460 26229
rect 17388 26139 17407 26173
rect 17441 26139 17460 26173
rect 17388 26083 17460 26139
rect 17388 26049 17407 26083
rect 17441 26049 17460 26083
rect 17388 25993 17460 26049
rect 17388 25959 17407 25993
rect 17441 25959 17460 25993
rect 16498 25888 16517 25922
rect 16551 25888 16570 25922
rect 16498 25865 16570 25888
rect 17388 25903 17460 25959
rect 17388 25869 17407 25903
rect 17441 25869 17460 25903
rect 17388 25865 17460 25869
rect 16498 25846 17460 25865
rect 16498 25812 16575 25846
rect 16609 25812 16665 25846
rect 16699 25812 16755 25846
rect 16789 25812 16845 25846
rect 16879 25812 16935 25846
rect 16969 25812 17025 25846
rect 17059 25812 17115 25846
rect 17149 25812 17205 25846
rect 17239 25812 17295 25846
rect 17329 25812 17460 25846
rect 16498 25793 17460 25812
rect 13810 25392 14772 25411
rect 13810 25358 13921 25392
rect 13955 25358 14011 25392
rect 14045 25358 14101 25392
rect 14135 25358 14191 25392
rect 14225 25358 14281 25392
rect 14315 25358 14371 25392
rect 14405 25358 14461 25392
rect 14495 25358 14551 25392
rect 14585 25358 14641 25392
rect 14675 25358 14772 25392
rect 13810 25339 14772 25358
rect 13810 25298 13882 25339
rect 13810 25264 13829 25298
rect 13863 25264 13882 25298
rect 14700 25279 14772 25339
rect 13810 25208 13882 25264
rect 13810 25174 13829 25208
rect 13863 25174 13882 25208
rect 13810 25118 13882 25174
rect 13810 25084 13829 25118
rect 13863 25084 13882 25118
rect 13810 25028 13882 25084
rect 13810 24994 13829 25028
rect 13863 24994 13882 25028
rect 13810 24938 13882 24994
rect 13810 24904 13829 24938
rect 13863 24904 13882 24938
rect 13810 24848 13882 24904
rect 13810 24814 13829 24848
rect 13863 24814 13882 24848
rect 13810 24758 13882 24814
rect 13810 24724 13829 24758
rect 13863 24724 13882 24758
rect 13810 24668 13882 24724
rect 13810 24634 13829 24668
rect 13863 24634 13882 24668
rect 13810 24578 13882 24634
rect 14700 25245 14719 25279
rect 14753 25245 14772 25279
rect 14700 25189 14772 25245
rect 14700 25155 14719 25189
rect 14753 25155 14772 25189
rect 14700 25099 14772 25155
rect 14700 25065 14719 25099
rect 14753 25065 14772 25099
rect 14700 25009 14772 25065
rect 14700 24975 14719 25009
rect 14753 24975 14772 25009
rect 14700 24919 14772 24975
rect 14700 24885 14719 24919
rect 14753 24885 14772 24919
rect 14700 24829 14772 24885
rect 14700 24795 14719 24829
rect 14753 24795 14772 24829
rect 14700 24739 14772 24795
rect 14700 24705 14719 24739
rect 14753 24705 14772 24739
rect 14700 24649 14772 24705
rect 14700 24615 14719 24649
rect 14753 24615 14772 24649
rect 13810 24544 13829 24578
rect 13863 24544 13882 24578
rect 13810 24521 13882 24544
rect 14700 24559 14772 24615
rect 14700 24525 14719 24559
rect 14753 24525 14772 24559
rect 14700 24521 14772 24525
rect 13810 24502 14772 24521
rect 13810 24468 13887 24502
rect 13921 24468 13977 24502
rect 14011 24468 14067 24502
rect 14101 24468 14157 24502
rect 14191 24468 14247 24502
rect 14281 24468 14337 24502
rect 14371 24468 14427 24502
rect 14461 24468 14517 24502
rect 14551 24468 14607 24502
rect 14641 24468 14772 24502
rect 13810 24449 14772 24468
rect 15154 25392 16116 25411
rect 15154 25358 15265 25392
rect 15299 25358 15355 25392
rect 15389 25358 15445 25392
rect 15479 25358 15535 25392
rect 15569 25358 15625 25392
rect 15659 25358 15715 25392
rect 15749 25358 15805 25392
rect 15839 25358 15895 25392
rect 15929 25358 15985 25392
rect 16019 25358 16116 25392
rect 15154 25339 16116 25358
rect 15154 25298 15226 25339
rect 15154 25264 15173 25298
rect 15207 25264 15226 25298
rect 16044 25279 16116 25339
rect 15154 25208 15226 25264
rect 15154 25174 15173 25208
rect 15207 25174 15226 25208
rect 15154 25118 15226 25174
rect 15154 25084 15173 25118
rect 15207 25084 15226 25118
rect 15154 25028 15226 25084
rect 15154 24994 15173 25028
rect 15207 24994 15226 25028
rect 15154 24938 15226 24994
rect 15154 24904 15173 24938
rect 15207 24904 15226 24938
rect 15154 24848 15226 24904
rect 15154 24814 15173 24848
rect 15207 24814 15226 24848
rect 15154 24758 15226 24814
rect 15154 24724 15173 24758
rect 15207 24724 15226 24758
rect 15154 24668 15226 24724
rect 15154 24634 15173 24668
rect 15207 24634 15226 24668
rect 15154 24578 15226 24634
rect 16044 25245 16063 25279
rect 16097 25245 16116 25279
rect 16044 25189 16116 25245
rect 16044 25155 16063 25189
rect 16097 25155 16116 25189
rect 16044 25099 16116 25155
rect 16044 25065 16063 25099
rect 16097 25065 16116 25099
rect 16044 25009 16116 25065
rect 16044 24975 16063 25009
rect 16097 24975 16116 25009
rect 16044 24919 16116 24975
rect 16044 24885 16063 24919
rect 16097 24885 16116 24919
rect 16044 24829 16116 24885
rect 16044 24795 16063 24829
rect 16097 24795 16116 24829
rect 16044 24739 16116 24795
rect 16044 24705 16063 24739
rect 16097 24705 16116 24739
rect 16044 24649 16116 24705
rect 16044 24615 16063 24649
rect 16097 24615 16116 24649
rect 15154 24544 15173 24578
rect 15207 24544 15226 24578
rect 15154 24521 15226 24544
rect 16044 24559 16116 24615
rect 16044 24525 16063 24559
rect 16097 24525 16116 24559
rect 16044 24521 16116 24525
rect 15154 24502 16116 24521
rect 15154 24468 15231 24502
rect 15265 24468 15321 24502
rect 15355 24468 15411 24502
rect 15445 24468 15501 24502
rect 15535 24468 15591 24502
rect 15625 24468 15681 24502
rect 15715 24468 15771 24502
rect 15805 24468 15861 24502
rect 15895 24468 15951 24502
rect 15985 24468 16116 24502
rect 15154 24449 16116 24468
rect 16498 25392 17460 25411
rect 16498 25358 16609 25392
rect 16643 25358 16699 25392
rect 16733 25358 16789 25392
rect 16823 25358 16879 25392
rect 16913 25358 16969 25392
rect 17003 25358 17059 25392
rect 17093 25358 17149 25392
rect 17183 25358 17239 25392
rect 17273 25358 17329 25392
rect 17363 25358 17460 25392
rect 16498 25339 17460 25358
rect 16498 25298 16570 25339
rect 16498 25264 16517 25298
rect 16551 25264 16570 25298
rect 17388 25279 17460 25339
rect 16498 25208 16570 25264
rect 16498 25174 16517 25208
rect 16551 25174 16570 25208
rect 16498 25118 16570 25174
rect 16498 25084 16517 25118
rect 16551 25084 16570 25118
rect 16498 25028 16570 25084
rect 16498 24994 16517 25028
rect 16551 24994 16570 25028
rect 16498 24938 16570 24994
rect 16498 24904 16517 24938
rect 16551 24904 16570 24938
rect 16498 24848 16570 24904
rect 16498 24814 16517 24848
rect 16551 24814 16570 24848
rect 16498 24758 16570 24814
rect 16498 24724 16517 24758
rect 16551 24724 16570 24758
rect 16498 24668 16570 24724
rect 16498 24634 16517 24668
rect 16551 24634 16570 24668
rect 16498 24578 16570 24634
rect 17388 25245 17407 25279
rect 17441 25245 17460 25279
rect 17388 25189 17460 25245
rect 17388 25155 17407 25189
rect 17441 25155 17460 25189
rect 17388 25099 17460 25155
rect 17388 25065 17407 25099
rect 17441 25065 17460 25099
rect 17388 25009 17460 25065
rect 17388 24975 17407 25009
rect 17441 24975 17460 25009
rect 17388 24919 17460 24975
rect 17388 24885 17407 24919
rect 17441 24885 17460 24919
rect 17388 24829 17460 24885
rect 17388 24795 17407 24829
rect 17441 24795 17460 24829
rect 17388 24739 17460 24795
rect 17388 24705 17407 24739
rect 17441 24705 17460 24739
rect 17388 24649 17460 24705
rect 17388 24615 17407 24649
rect 17441 24615 17460 24649
rect 16498 24544 16517 24578
rect 16551 24544 16570 24578
rect 16498 24521 16570 24544
rect 17388 24559 17460 24615
rect 17388 24525 17407 24559
rect 17441 24525 17460 24559
rect 17388 24521 17460 24525
rect 16498 24502 17460 24521
rect 16498 24468 16575 24502
rect 16609 24468 16665 24502
rect 16699 24468 16755 24502
rect 16789 24468 16845 24502
rect 16879 24468 16935 24502
rect 16969 24468 17025 24502
rect 17059 24468 17115 24502
rect 17149 24468 17205 24502
rect 17239 24468 17295 24502
rect 17329 24468 17460 24502
rect 16498 24449 17460 24468
<< mvpsubdiff >>
rect 5930 24236 10848 24248
rect 5930 24202 6038 24236
rect 6366 24202 6524 24236
rect 6852 24202 7010 24236
rect 7338 24202 7496 24236
rect 7824 24202 7982 24236
rect 8310 24202 8468 24236
rect 8796 24202 8954 24236
rect 9282 24202 9440 24236
rect 9768 24202 9926 24236
rect 10254 24202 10412 24236
rect 10740 24202 10848 24236
rect 5930 24190 10848 24202
rect 5930 24140 5988 24190
rect 5930 19972 5942 24140
rect 5976 19972 5988 24140
rect 6416 24140 6474 24190
rect 5930 19922 5988 19972
rect 6416 19972 6428 24140
rect 6462 19972 6474 24140
rect 6902 24140 6960 24190
rect 6416 19922 6474 19972
rect 6902 19972 6914 24140
rect 6948 19972 6960 24140
rect 7388 24140 7446 24190
rect 6902 19922 6960 19972
rect 7388 19972 7400 24140
rect 7434 19972 7446 24140
rect 7874 24140 7932 24190
rect 7388 19922 7446 19972
rect 7874 19972 7886 24140
rect 7920 19972 7932 24140
rect 8360 24140 8418 24190
rect 7874 19922 7932 19972
rect 8360 19972 8372 24140
rect 8406 19972 8418 24140
rect 8846 24140 8904 24190
rect 8360 19922 8418 19972
rect 8846 19972 8858 24140
rect 8892 19972 8904 24140
rect 9332 24140 9390 24190
rect 8846 19922 8904 19972
rect 9332 19972 9344 24140
rect 9378 19972 9390 24140
rect 9818 24140 9876 24190
rect 9332 19922 9390 19972
rect 9818 19972 9830 24140
rect 9864 19972 9876 24140
rect 10304 24140 10362 24190
rect 9818 19922 9876 19972
rect 10304 19972 10316 24140
rect 10350 19972 10362 24140
rect 10790 24140 10848 24190
rect 10304 19922 10362 19972
rect 10790 19972 10802 24140
rect 10836 19972 10848 24140
rect 15651 23829 20035 23841
rect 15651 23795 15759 23829
rect 19927 23795 20035 23829
rect 15651 23783 20035 23795
rect 15651 23733 15709 23783
rect 11195 23429 15579 23441
rect 11195 23395 11303 23429
rect 15471 23395 15579 23429
rect 11195 23383 15579 23395
rect 11195 23333 11253 23383
rect 11195 22505 11207 23333
rect 11241 22505 11253 23333
rect 15521 23333 15579 23383
rect 11195 22455 11253 22505
rect 15521 22505 15533 23333
rect 15567 22505 15579 23333
rect 15521 22455 15579 22505
rect 11195 22443 15579 22455
rect 11195 22409 11303 22443
rect 15471 22409 15579 22443
rect 11195 22397 15579 22409
rect 15651 22505 15663 23733
rect 15697 22505 15709 23733
rect 19977 23733 20035 23783
rect 15651 22455 15709 22505
rect 19977 22505 19989 23733
rect 20023 22505 20035 23733
rect 19977 22455 20035 22505
rect 15651 22443 20035 22455
rect 15651 22409 15759 22443
rect 19927 22409 20035 22443
rect 15651 22397 20035 22409
rect 11202 22157 15586 22169
rect 11202 22123 11310 22157
rect 15478 22123 15586 22157
rect 11202 22111 15586 22123
rect 11202 22061 11260 22111
rect 11202 20833 11214 22061
rect 11248 20833 11260 22061
rect 15528 22061 15586 22111
rect 11202 20783 11260 20833
rect 15528 20833 15540 22061
rect 15574 20833 15586 22061
rect 15651 22157 20035 22169
rect 15651 22123 15759 22157
rect 19927 22123 20035 22157
rect 15651 22111 20035 22123
rect 15651 22061 15709 22111
rect 15651 21233 15663 22061
rect 15697 21233 15709 22061
rect 19977 22061 20035 22111
rect 15651 21183 15709 21233
rect 19977 21233 19989 22061
rect 20023 21233 20035 22061
rect 19977 21183 20035 21233
rect 15651 21171 20035 21183
rect 15651 21137 15759 21171
rect 19927 21137 20035 21171
rect 15651 21125 20035 21137
rect 15528 20783 15586 20833
rect 11202 20771 15586 20783
rect 11202 20737 11310 20771
rect 15478 20737 15586 20771
rect 11202 20725 15586 20737
rect 10790 19922 10848 19972
rect 5930 19910 10848 19922
rect 5930 19876 6038 19910
rect 6366 19876 6524 19910
rect 6852 19876 7010 19910
rect 7338 19876 7496 19910
rect 7824 19876 7982 19910
rect 8310 19876 8468 19910
rect 8796 19876 8954 19910
rect 9282 19876 9440 19910
rect 9768 19876 9926 19910
rect 10254 19876 10412 19910
rect 10740 19876 10848 19910
rect 5930 19864 10848 19876
rect 11271 9860 11755 9872
rect 11271 9826 11379 9860
rect 11647 9826 11755 9860
rect 11271 9814 11755 9826
rect 11271 9764 11329 9814
rect 11271 9336 11283 9764
rect 11317 9336 11329 9764
rect 11697 9764 11755 9814
rect 11271 9286 11329 9336
rect 11697 9336 11709 9764
rect 11743 9336 11755 9764
rect 11697 9286 11755 9336
rect 11271 9274 11755 9286
rect 11271 9240 11379 9274
rect 11647 9240 11755 9274
rect 11271 9228 11755 9240
rect 11827 9860 12311 9872
rect 11827 9826 11935 9860
rect 12203 9826 12311 9860
rect 11827 9814 12311 9826
rect 11827 9764 11885 9814
rect 11827 9336 11839 9764
rect 11873 9336 11885 9764
rect 12253 9764 12311 9814
rect 11827 9286 11885 9336
rect 12253 9336 12265 9764
rect 12299 9336 12311 9764
rect 12253 9286 12311 9336
rect 11827 9274 12311 9286
rect 11827 9240 11935 9274
rect 12203 9240 12311 9274
rect 11827 9228 12311 9240
rect 12383 9860 12867 9872
rect 12383 9826 12491 9860
rect 12759 9826 12867 9860
rect 12383 9814 12867 9826
rect 12383 9764 12441 9814
rect 12383 9336 12395 9764
rect 12429 9336 12441 9764
rect 12809 9764 12867 9814
rect 12383 9286 12441 9336
rect 12809 9336 12821 9764
rect 12855 9336 12867 9764
rect 12809 9286 12867 9336
rect 12383 9274 12867 9286
rect 12383 9240 12491 9274
rect 12759 9240 12867 9274
rect 12383 9228 12867 9240
rect 12939 9860 13423 9872
rect 12939 9826 13047 9860
rect 13315 9826 13423 9860
rect 12939 9814 13423 9826
rect 12939 9764 12997 9814
rect 12939 9336 12951 9764
rect 12985 9336 12997 9764
rect 13365 9764 13423 9814
rect 12939 9286 12997 9336
rect 13365 9336 13377 9764
rect 13411 9336 13423 9764
rect 13365 9286 13423 9336
rect 12939 9274 13423 9286
rect 12939 9240 13047 9274
rect 13315 9240 13423 9274
rect 12939 9228 13423 9240
rect 5319 8609 6903 8621
rect 5319 8575 5427 8609
rect 6795 8575 6903 8609
rect 5319 8563 6903 8575
rect 5319 8513 5377 8563
rect 5319 8085 5331 8513
rect 5365 8085 5377 8513
rect 6845 8513 6903 8563
rect 5319 8035 5377 8085
rect 6845 8085 6857 8513
rect 6891 8085 6903 8513
rect 6845 8035 6903 8085
rect 5319 8023 6903 8035
rect 5319 7989 5427 8023
rect 6795 7989 6903 8023
rect 5319 7977 6903 7989
rect 6975 8609 8559 8621
rect 6975 8575 7083 8609
rect 8451 8575 8559 8609
rect 6975 8563 8559 8575
rect 6975 8513 7033 8563
rect 6975 8085 6987 8513
rect 7021 8085 7033 8513
rect 8501 8513 8559 8563
rect 6975 8035 7033 8085
rect 8501 8085 8513 8513
rect 8547 8085 8559 8513
rect 8501 8035 8559 8085
rect 6975 8023 8559 8035
rect 6975 7989 7083 8023
rect 8451 7989 8559 8023
rect 6975 7977 8559 7989
rect 8905 8609 9729 8621
rect 8905 8575 9013 8609
rect 9621 8575 9729 8609
rect 8905 8563 9729 8575
rect 8905 8513 8963 8563
rect 8905 8085 8917 8513
rect 8951 8085 8963 8513
rect 9671 8513 9729 8563
rect 8905 8035 8963 8085
rect 9671 8085 9683 8513
rect 9717 8085 9729 8513
rect 9671 8035 9729 8085
rect 8905 8023 9729 8035
rect 8905 7989 9013 8023
rect 9621 7989 9729 8023
rect 8905 7977 9729 7989
rect 9877 8610 10701 8622
rect 9877 8576 9985 8610
rect 10593 8576 10701 8610
rect 9877 8564 10701 8576
rect 9877 8514 9935 8564
rect 9877 8086 9889 8514
rect 9923 8086 9935 8514
rect 10643 8514 10701 8564
rect 9877 8036 9935 8086
rect 10643 8086 10655 8514
rect 10689 8086 10701 8514
rect 10643 8036 10701 8086
rect 9877 8024 10701 8036
rect 9877 7990 9985 8024
rect 10593 7990 10701 8024
rect 9877 7978 10701 7990
rect 5319 7893 6903 7905
rect 5319 7859 5427 7893
rect 6795 7859 6903 7893
rect 5319 7847 6903 7859
rect 5319 7797 5377 7847
rect 5319 7369 5331 7797
rect 5365 7369 5377 7797
rect 6845 7797 6903 7847
rect 5319 7319 5377 7369
rect 6845 7369 6857 7797
rect 6891 7369 6903 7797
rect 6845 7319 6903 7369
rect 5319 7307 6903 7319
rect 5319 7273 5427 7307
rect 6795 7273 6903 7307
rect 5319 7261 6903 7273
rect 6975 7893 8559 7905
rect 6975 7859 7083 7893
rect 8451 7859 8559 7893
rect 6975 7847 8559 7859
rect 6975 7797 7033 7847
rect 6975 7369 6987 7797
rect 7021 7369 7033 7797
rect 8501 7797 8559 7847
rect 6975 7319 7033 7369
rect 8501 7369 8513 7797
rect 8547 7369 8559 7797
rect 8501 7319 8559 7369
rect 6975 7307 8559 7319
rect 6975 7273 7083 7307
rect 8451 7273 8559 7307
rect 6975 7261 8559 7273
rect 5319 7177 6903 7189
rect 5319 7143 5427 7177
rect 6795 7143 6903 7177
rect 5319 7131 6903 7143
rect 5319 7081 5377 7131
rect 5319 6653 5331 7081
rect 5365 6653 5377 7081
rect 6845 7081 6903 7131
rect 5319 6603 5377 6653
rect 6845 6653 6857 7081
rect 6891 6653 6903 7081
rect 6845 6603 6903 6653
rect 5319 6591 6903 6603
rect 5319 6557 5427 6591
rect 6795 6557 6903 6591
rect 5319 6545 6903 6557
rect 6975 7177 8559 7189
rect 6975 7143 7083 7177
rect 8451 7143 8559 7177
rect 6975 7131 8559 7143
rect 6975 7081 7033 7131
rect 6975 6653 6987 7081
rect 7021 6653 7033 7081
rect 8501 7081 8559 7131
rect 6975 6603 7033 6653
rect 8501 6653 8513 7081
rect 8547 6653 8559 7081
rect 8501 6603 8559 6653
rect 6975 6591 8559 6603
rect 6975 6557 7083 6591
rect 8451 6557 8559 6591
rect 6975 6545 8559 6557
rect 16463 9898 20265 9910
rect 16463 9864 16571 9898
rect 20157 9864 20265 9898
rect 16463 9852 20265 9864
rect 16463 9802 16521 9852
rect 16463 7574 16475 9802
rect 16509 7574 16521 9802
rect 20207 9802 20265 9852
rect 16463 7524 16521 7574
rect 20207 7574 20219 9802
rect 20253 7574 20265 9802
rect 20207 7524 20265 7574
rect 16463 7512 20265 7524
rect 16463 7478 16571 7512
rect 20157 7478 20265 7512
rect 16463 7466 20265 7478
rect 21515 8079 23959 8091
rect 21515 8045 21623 8079
rect 23851 8045 23959 8079
rect 21515 8033 23959 8045
rect 21515 7983 21573 8033
rect 5319 6461 6903 6473
rect 5319 6427 5427 6461
rect 6795 6427 6903 6461
rect 5319 6415 6903 6427
rect 5319 6365 5377 6415
rect 5319 5937 5331 6365
rect 5365 5937 5377 6365
rect 6845 6365 6903 6415
rect 5319 5887 5377 5937
rect 6845 5937 6857 6365
rect 6891 5937 6903 6365
rect 6845 5887 6903 5937
rect 5319 5875 6903 5887
rect 5319 5841 5427 5875
rect 6795 5841 6903 5875
rect 5319 5829 6903 5841
rect 6975 6461 8559 6473
rect 6975 6427 7083 6461
rect 8451 6427 8559 6461
rect 6975 6415 8559 6427
rect 6975 6365 7033 6415
rect 6975 5937 6987 6365
rect 7021 5937 7033 6365
rect 8501 6365 8559 6415
rect 6975 5887 7033 5937
rect 8501 5937 8513 6365
rect 8547 5937 8559 6365
rect 8501 5887 8559 5937
rect 6975 5875 8559 5887
rect 6975 5841 7083 5875
rect 8451 5841 8559 5875
rect 6975 5829 8559 5841
rect 16459 7311 18275 7323
rect 16459 7277 16567 7311
rect 16995 7277 17153 7311
rect 17581 7277 17739 7311
rect 18167 7277 18275 7311
rect 16459 7265 18275 7277
rect 16459 7215 16517 7265
rect 16459 5047 16471 7215
rect 16505 5047 16517 7215
rect 17045 7215 17103 7265
rect 16459 4997 16517 5047
rect 17045 5047 17057 7215
rect 17091 5047 17103 7215
rect 17631 7215 17689 7265
rect 17045 4997 17103 5047
rect 17631 5047 17643 7215
rect 17677 5047 17689 7215
rect 18217 7215 18275 7265
rect 17631 4997 17689 5047
rect 18217 5047 18229 7215
rect 18263 5047 18275 7215
rect 18217 4997 18275 5047
rect 16459 4985 18275 4997
rect 16459 4951 16567 4985
rect 16995 4951 17153 4985
rect 17581 4951 17739 4985
rect 18167 4951 18275 4985
rect 16459 4939 18275 4951
rect 16459 4849 18275 4861
rect 16459 4815 16567 4849
rect 16995 4815 17153 4849
rect 17581 4815 17739 4849
rect 18167 4815 18275 4849
rect 16459 4803 18275 4815
rect 16459 4753 16517 4803
rect 16459 2585 16471 4753
rect 16505 2585 16517 4753
rect 17045 4753 17103 4803
rect 16459 2535 16517 2585
rect 17045 2585 17057 4753
rect 17091 2585 17103 4753
rect 17631 4753 17689 4803
rect 17045 2535 17103 2585
rect 17631 2585 17643 4753
rect 17677 2585 17689 4753
rect 18217 4753 18275 4803
rect 17631 2535 17689 2585
rect 18217 2585 18229 4753
rect 18263 2585 18275 4753
rect 18217 2535 18275 2585
rect 16459 2523 18275 2535
rect 16459 2489 16567 2523
rect 16995 2489 17153 2523
rect 17581 2489 17739 2523
rect 18167 2489 18275 2523
rect 16459 2477 18275 2489
rect 21515 6015 21527 7983
rect 21561 6015 21573 7983
rect 23901 7983 23959 8033
rect 21515 5965 21573 6015
rect 23901 6015 23913 7983
rect 23947 6015 23959 7983
rect 23901 5965 23959 6015
rect 21515 5953 23959 5965
rect 21515 5919 21623 5953
rect 23851 5919 23959 5953
rect 21515 5907 23959 5919
rect 21515 5829 23959 5841
rect 21515 5795 21623 5829
rect 23851 5795 23959 5829
rect 21515 5783 23959 5795
rect 21515 5733 21573 5783
rect 21515 3765 21527 5733
rect 21561 3765 21573 5733
rect 23901 5733 23959 5783
rect 21515 3715 21573 3765
rect 23901 3765 23913 5733
rect 23947 3765 23959 5733
rect 23901 3715 23959 3765
rect 21515 3703 23959 3715
rect 21515 3669 21623 3703
rect 23851 3669 23959 3703
rect 21515 3657 23959 3669
rect 24444 3971 26888 3983
rect 24444 3937 24552 3971
rect 26780 3937 26888 3971
rect 24444 3925 26888 3937
rect 24444 3875 24502 3925
rect 21300 3137 24206 3149
rect 21300 3103 21408 3137
rect 24098 3103 24206 3137
rect 21300 3091 24206 3103
rect 21300 3041 21358 3091
rect 21300 1813 21312 3041
rect 21346 1813 21358 3041
rect 24148 3041 24206 3091
rect 21300 1763 21358 1813
rect 24148 1813 24160 3041
rect 24194 1813 24206 3041
rect 24148 1763 24206 1813
rect 24444 1907 24456 3875
rect 24490 1907 24502 3875
rect 26830 3875 26888 3925
rect 24444 1857 24502 1907
rect 26830 1907 26842 3875
rect 26876 1907 26888 3875
rect 26830 1857 26888 1907
rect 24444 1845 26888 1857
rect 24444 1811 24552 1845
rect 26780 1811 26888 1845
rect 24444 1799 26888 1811
rect 21300 1751 24206 1763
rect 21300 1717 21408 1751
rect 24098 1717 24206 1751
rect 21300 1705 24206 1717
<< mvnsubdiff >>
rect 6087 31137 10797 31149
rect 6087 31103 6195 31137
rect 8363 31103 8521 31137
rect 10689 31103 10797 31137
rect 6087 31091 10797 31103
rect 6087 31041 6145 31091
rect 6087 30595 6099 31041
rect 6133 30595 6145 31041
rect 8413 31041 8471 31091
rect 6087 30545 6145 30595
rect 8413 30595 8425 31041
rect 8459 30595 8471 31041
rect 10739 31041 10797 31091
rect 8413 30545 8471 30595
rect 10739 30595 10751 31041
rect 10785 30595 10797 31041
rect 10739 30545 10797 30595
rect 6087 30533 10797 30545
rect 6087 30499 6195 30533
rect 8363 30499 8521 30533
rect 10689 30499 10797 30533
rect 6087 30487 10797 30499
rect 6212 19270 10596 19282
rect 6212 19236 6320 19270
rect 10488 19236 10596 19270
rect 6212 19224 10596 19236
rect 6212 19174 6270 19224
rect 6212 18092 6224 19174
rect 6258 18092 6270 19174
rect 10538 19174 10596 19224
rect 6212 18042 6270 18092
rect 10538 18092 10550 19174
rect 10584 18092 10596 19174
rect 10538 18042 10596 18092
rect 6212 18030 10596 18042
rect 6212 17996 6320 18030
rect 10488 17996 10596 18030
rect 6212 17984 10596 17996
rect 11300 19270 20010 19282
rect 11300 19236 11408 19270
rect 15576 19236 15734 19270
rect 19902 19236 20010 19270
rect 11300 19224 20010 19236
rect 11300 19174 11358 19224
rect 6212 17870 10596 17882
rect 6212 17836 6320 17870
rect 10488 17836 10596 17870
rect 6212 17824 10596 17836
rect 6212 17774 6270 17824
rect 6212 16928 6224 17774
rect 6258 16928 6270 17774
rect 10538 17774 10596 17824
rect 6212 16878 6270 16928
rect 10538 16928 10550 17774
rect 10584 16928 10596 17774
rect 10538 16878 10596 16928
rect 6212 16866 10596 16878
rect 6212 16832 6320 16866
rect 10488 16832 10596 16866
rect 6212 16820 10596 16832
rect 11300 16928 11312 19174
rect 11346 16928 11358 19174
rect 15626 19174 15684 19224
rect 11300 16878 11358 16928
rect 15626 16928 15638 19174
rect 15672 16928 15684 19174
rect 19952 19174 20010 19224
rect 15626 16878 15684 16928
rect 19952 16928 19964 19174
rect 19998 16928 20010 19174
rect 19952 16878 20010 16928
rect 11300 16866 20010 16878
rect 11300 16832 11408 16866
rect 15576 16832 15734 16866
rect 19902 16832 20010 16866
rect 11300 16820 20010 16832
rect 11300 16770 11358 16820
rect 8222 15066 10596 15078
rect 8222 15032 8330 15066
rect 10488 15032 10596 15066
rect 8222 15020 10596 15032
rect 8222 14970 8280 15020
rect 8222 14524 8234 14970
rect 8268 14524 8280 14970
rect 10538 14970 10596 15020
rect 8222 14474 8280 14524
rect 10538 14524 10550 14970
rect 10584 14524 10596 14970
rect 10538 14474 10596 14524
rect 8222 14462 10596 14474
rect 8222 14428 8330 14462
rect 10488 14428 10596 14462
rect 8222 14416 10596 14428
rect 11300 14524 11312 16770
rect 11346 14524 11358 16770
rect 15626 16770 15684 16820
rect 11300 14474 11358 14524
rect 15626 14524 15638 16770
rect 15672 14524 15684 16770
rect 19952 16770 20010 16820
rect 15626 14474 15684 14524
rect 19952 14524 19964 16770
rect 19998 14524 20010 16770
rect 20668 18902 21734 18914
rect 20668 18868 20776 18902
rect 21122 18868 21280 18902
rect 21626 18868 21734 18902
rect 20668 18856 21734 18868
rect 20668 18806 20726 18856
rect 20668 14638 20680 18806
rect 20714 14638 20726 18806
rect 21172 18806 21230 18856
rect 20668 14588 20726 14638
rect 21172 14638 21184 18806
rect 21218 14638 21230 18806
rect 21676 18806 21734 18856
rect 21172 14588 21230 14638
rect 21676 14638 21688 18806
rect 21722 14638 21734 18806
rect 21676 14588 21734 14638
rect 20668 14576 21734 14588
rect 20668 14542 20776 14576
rect 21122 14542 21280 14576
rect 21626 14542 21734 14576
rect 20668 14530 21734 14542
rect 19952 14474 20010 14524
rect 11300 14462 20010 14474
rect 11300 14428 11408 14462
rect 15576 14428 15734 14462
rect 19902 14428 20010 14462
rect 11300 14416 20010 14428
rect 7927 12542 10321 12554
rect 7927 12508 8035 12542
rect 10213 12508 10321 12542
rect 7927 12496 10321 12508
rect 7927 12446 7985 12496
rect 7927 12000 7939 12446
rect 7973 12000 7985 12446
rect 10263 12446 10321 12496
rect 7927 11950 7985 12000
rect 10263 12000 10275 12446
rect 10309 12000 10321 12446
rect 10263 11950 10321 12000
rect 7927 11938 10321 11950
rect 7927 11904 8035 11938
rect 10213 11904 10321 11938
rect 7927 11892 10321 11904
rect 5927 11779 10311 11791
rect 5927 11745 6035 11779
rect 10203 11745 10311 11779
rect 5927 11733 10311 11745
rect 5927 11683 5985 11733
rect 5927 11037 5939 11683
rect 5973 11037 5985 11683
rect 10253 11683 10311 11733
rect 5927 10987 5985 11037
rect 10253 11037 10265 11683
rect 10299 11037 10311 11683
rect 10253 10987 10311 11037
rect 5927 10975 10311 10987
rect 5927 10941 6035 10975
rect 10203 10941 10311 10975
rect 5927 10929 10311 10941
rect 11913 11015 11973 11049
rect 12757 11015 12817 11049
rect 11913 10989 11947 11015
rect 8905 10811 9769 10823
rect 6039 10793 6903 10805
rect 6039 10759 6147 10793
rect 6795 10759 6903 10793
rect 6039 10747 6903 10759
rect 6039 10697 6097 10747
rect 6039 9951 6051 10697
rect 6085 9951 6097 10697
rect 6845 10697 6903 10747
rect 6039 9901 6097 9951
rect 6845 9951 6857 10697
rect 6891 9951 6903 10697
rect 6845 9901 6903 9951
rect 6039 9889 6903 9901
rect 6039 9855 6147 9889
rect 6795 9855 6903 9889
rect 6039 9843 6903 9855
rect 6975 10793 7839 10805
rect 6975 10759 7083 10793
rect 7731 10759 7839 10793
rect 6975 10747 7839 10759
rect 6975 10697 7033 10747
rect 6975 9951 6987 10697
rect 7021 9951 7033 10697
rect 7781 10697 7839 10747
rect 6975 9901 7033 9951
rect 7781 9951 7793 10697
rect 7827 9951 7839 10697
rect 7781 9901 7839 9951
rect 6975 9889 7839 9901
rect 6975 9855 7083 9889
rect 7731 9855 7839 9889
rect 8905 10777 9013 10811
rect 9661 10777 9769 10811
rect 8905 10765 9769 10777
rect 8905 10715 8963 10765
rect 8905 9969 8917 10715
rect 8951 9969 8963 10715
rect 9711 10715 9769 10765
rect 8905 9919 8963 9969
rect 9711 9969 9723 10715
rect 9757 9969 9769 10715
rect 9711 9919 9769 9969
rect 8905 9907 9769 9919
rect 8905 9873 9013 9907
rect 9661 9873 9769 9907
rect 8905 9861 9769 9873
rect 9837 10811 10701 10823
rect 9837 10777 9945 10811
rect 10593 10777 10701 10811
rect 9837 10765 10701 10777
rect 9837 10715 9895 10765
rect 9837 9969 9849 10715
rect 9883 9969 9895 10715
rect 10643 10715 10701 10765
rect 9837 9919 9895 9969
rect 10643 9969 10655 10715
rect 10689 9969 10701 10715
rect 12783 10989 12817 11015
rect 11913 10507 11947 10533
rect 12783 10507 12817 10533
rect 11913 10473 11973 10507
rect 12757 10473 12817 10507
rect 10643 9919 10701 9969
rect 9837 9907 10701 9919
rect 9837 9873 9945 9907
rect 10593 9873 10701 9907
rect 9837 9861 10701 9873
rect 6975 9843 7839 9855
rect 6039 9751 6903 9763
rect 6039 9717 6147 9751
rect 6795 9717 6903 9751
rect 6039 9705 6903 9717
rect 6039 9655 6097 9705
rect 6039 8909 6051 9655
rect 6085 8909 6097 9655
rect 6845 9655 6903 9705
rect 6039 8859 6097 8909
rect 6845 8909 6857 9655
rect 6891 8909 6903 9655
rect 6845 8859 6903 8909
rect 6039 8847 6903 8859
rect 6039 8813 6147 8847
rect 6795 8813 6903 8847
rect 6039 8801 6903 8813
rect 6975 9751 7839 9763
rect 6975 9717 7083 9751
rect 7731 9717 7839 9751
rect 6975 9705 7839 9717
rect 6975 9655 7033 9705
rect 6975 8909 6987 9655
rect 7021 8909 7033 9655
rect 7781 9655 7839 9705
rect 6975 8859 7033 8909
rect 7781 8909 7793 9655
rect 7827 8909 7839 9655
rect 7781 8859 7839 8909
rect 6975 8847 7839 8859
rect 6975 8813 7083 8847
rect 7731 8813 7839 8847
rect 6975 8801 7839 8813
rect 8905 9726 9769 9738
rect 8905 9692 9013 9726
rect 9661 9692 9769 9726
rect 8905 9680 9769 9692
rect 8905 9630 8963 9680
rect 8905 8884 8917 9630
rect 8951 8884 8963 9630
rect 9711 9630 9769 9680
rect 8905 8834 8963 8884
rect 9711 8884 9723 9630
rect 9757 8884 9769 9630
rect 9711 8834 9769 8884
rect 8905 8822 9769 8834
rect 8905 8788 9013 8822
rect 9661 8788 9769 8822
rect 8905 8776 9769 8788
rect 9837 9726 10701 9738
rect 9837 9692 9945 9726
rect 10593 9692 10701 9726
rect 9837 9680 10701 9692
rect 9837 9630 9895 9680
rect 9837 8884 9849 9630
rect 9883 8884 9895 9630
rect 10643 9630 10701 9680
rect 9837 8834 9895 8884
rect 10643 8884 10655 9630
rect 10689 8884 10701 9630
rect 10643 8834 10701 8884
rect 9837 8822 10701 8834
rect 9837 8788 9945 8822
rect 10593 8788 10701 8822
rect 9837 8776 10701 8788
rect 24600 8079 25862 8091
rect 24600 8045 24708 8079
rect 25754 8045 25862 8079
rect 24600 8033 25862 8045
rect 24600 7983 24658 8033
rect 24600 7615 24612 7983
rect 24646 7615 24658 7983
rect 25804 7983 25862 8033
rect 24600 7565 24658 7615
rect 25804 7615 25816 7983
rect 25850 7615 25862 7983
rect 25804 7565 25862 7615
rect 24600 7553 25862 7565
rect 24600 7519 24708 7553
rect 25754 7519 25862 7553
rect 24600 7507 25862 7519
rect 24600 7373 26762 7385
rect 24600 7339 24708 7373
rect 26654 7339 26762 7373
rect 24600 7327 26762 7339
rect 24600 7277 24658 7327
rect 24600 5103 24612 7277
rect 24646 5103 24658 7277
rect 26704 7277 26762 7327
rect 24600 5053 24658 5103
rect 26704 5103 26716 7277
rect 26750 5103 26762 7277
rect 26704 5053 26762 5103
rect 24600 5041 26762 5053
rect 24600 5007 24708 5041
rect 26654 5007 26762 5041
rect 24600 4995 26762 5007
<< psubdiffcont >>
rect 2752 42334 2890 42368
rect 3048 42334 3186 42368
rect 3344 42334 3482 42368
rect 3640 42334 3778 42368
rect 3936 42334 4074 42368
rect 4232 42334 4370 42368
rect 4528 42334 4666 42368
rect 4824 42334 4962 42368
rect 5120 42334 5258 42368
rect 5416 42334 5554 42368
rect 2656 36372 2690 42272
rect 2952 36372 2986 42272
rect 3248 36372 3282 42272
rect 3544 36372 3578 42272
rect 3840 36372 3874 42272
rect 4136 36372 4170 42272
rect 4432 36372 4466 42272
rect 4728 36372 4762 42272
rect 5024 36372 5058 42272
rect 5320 36372 5354 42272
rect 5616 36372 5650 42272
rect 2752 36276 2890 36310
rect 3048 36276 3186 36310
rect 3344 36276 3482 36310
rect 3640 36276 3778 36310
rect 3936 36276 4074 36310
rect 4232 36276 4370 36310
rect 4528 36276 4666 36310
rect 4824 36276 4962 36310
rect 5120 36276 5258 36310
rect 5416 36276 5554 36310
rect 2656 30314 2690 36214
rect 2952 30314 2986 36214
rect 3248 30314 3282 36214
rect 3544 30314 3578 36214
rect 3840 30314 3874 36214
rect 4136 30314 4170 36214
rect 4432 30314 4466 36214
rect 4728 30314 4762 36214
rect 5024 30314 5058 36214
rect 5320 30314 5354 36214
rect 5616 30314 5650 36214
rect 2752 30218 2890 30252
rect 3048 30218 3186 30252
rect 3344 30218 3482 30252
rect 3640 30218 3778 30252
rect 3936 30218 4074 30252
rect 4232 30218 4370 30252
rect 4528 30218 4666 30252
rect 4824 30218 4962 30252
rect 5120 30218 5258 30252
rect 5416 30218 5554 30252
rect 7552 28209 10352 28243
rect 10510 28209 13310 28243
rect 7456 28009 7490 28147
rect 10414 28009 10448 28147
rect 13372 28009 13406 28147
rect 7552 27913 10352 27947
rect 10510 27913 13310 27947
rect 7456 27713 7490 27851
rect 10414 27713 10448 27851
rect 13372 27713 13406 27851
rect 7552 27617 10352 27651
rect 10510 27617 13310 27651
rect 7456 27417 7490 27555
rect 10414 27417 10448 27555
rect 13372 27417 13406 27555
rect 7552 27321 10352 27355
rect 10510 27321 13310 27355
rect 7456 27121 7490 27259
rect 10414 27121 10448 27259
rect 13372 27121 13406 27259
rect 7552 27025 10352 27059
rect 10510 27025 13310 27059
rect 7456 26825 7490 26963
rect 10414 26825 10448 26963
rect 13781 28196 13815 28230
rect 13871 28196 13905 28230
rect 13961 28196 13995 28230
rect 14051 28196 14085 28230
rect 14141 28196 14175 28230
rect 14231 28196 14265 28230
rect 14321 28196 14355 28230
rect 14411 28196 14445 28230
rect 14501 28196 14535 28230
rect 14591 28196 14625 28230
rect 14681 28196 14715 28230
rect 14771 28196 14805 28230
rect 13680 28112 13714 28146
rect 14867 28112 14901 28146
rect 13680 28022 13714 28056
rect 13680 27932 13714 27966
rect 13680 27842 13714 27876
rect 13680 27752 13714 27786
rect 13680 27662 13714 27696
rect 13680 27572 13714 27606
rect 13680 27482 13714 27516
rect 13680 27392 13714 27426
rect 13680 27302 13714 27336
rect 13680 27212 13714 27246
rect 13680 27122 13714 27156
rect 14867 28022 14901 28056
rect 14867 27932 14901 27966
rect 14867 27842 14901 27876
rect 14867 27752 14901 27786
rect 14867 27662 14901 27696
rect 14867 27572 14901 27606
rect 14867 27482 14901 27516
rect 14867 27392 14901 27426
rect 14867 27302 14901 27336
rect 14867 27212 14901 27246
rect 14867 27122 14901 27156
rect 13680 27032 13714 27066
rect 13781 27009 13815 27043
rect 13871 27009 13905 27043
rect 13961 27009 13995 27043
rect 14051 27009 14085 27043
rect 14141 27009 14175 27043
rect 14231 27009 14265 27043
rect 14321 27009 14355 27043
rect 14411 27009 14445 27043
rect 14501 27009 14535 27043
rect 14591 27009 14625 27043
rect 14681 27009 14715 27043
rect 14771 27009 14805 27043
rect 14867 27032 14901 27066
rect 15125 28196 15159 28230
rect 15215 28196 15249 28230
rect 15305 28196 15339 28230
rect 15395 28196 15429 28230
rect 15485 28196 15519 28230
rect 15575 28196 15609 28230
rect 15665 28196 15699 28230
rect 15755 28196 15789 28230
rect 15845 28196 15879 28230
rect 15935 28196 15969 28230
rect 16025 28196 16059 28230
rect 16115 28196 16149 28230
rect 15024 28112 15058 28146
rect 16211 28112 16245 28146
rect 15024 28022 15058 28056
rect 15024 27932 15058 27966
rect 15024 27842 15058 27876
rect 15024 27752 15058 27786
rect 15024 27662 15058 27696
rect 15024 27572 15058 27606
rect 15024 27482 15058 27516
rect 15024 27392 15058 27426
rect 15024 27302 15058 27336
rect 15024 27212 15058 27246
rect 15024 27122 15058 27156
rect 16211 28022 16245 28056
rect 16211 27932 16245 27966
rect 16211 27842 16245 27876
rect 16211 27752 16245 27786
rect 16211 27662 16245 27696
rect 16211 27572 16245 27606
rect 16211 27482 16245 27516
rect 16211 27392 16245 27426
rect 16211 27302 16245 27336
rect 16211 27212 16245 27246
rect 16211 27122 16245 27156
rect 15024 27032 15058 27066
rect 15125 27009 15159 27043
rect 15215 27009 15249 27043
rect 15305 27009 15339 27043
rect 15395 27009 15429 27043
rect 15485 27009 15519 27043
rect 15575 27009 15609 27043
rect 15665 27009 15699 27043
rect 15755 27009 15789 27043
rect 15845 27009 15879 27043
rect 15935 27009 15969 27043
rect 16025 27009 16059 27043
rect 16115 27009 16149 27043
rect 16211 27032 16245 27066
rect 16469 28196 16503 28230
rect 16559 28196 16593 28230
rect 16649 28196 16683 28230
rect 16739 28196 16773 28230
rect 16829 28196 16863 28230
rect 16919 28196 16953 28230
rect 17009 28196 17043 28230
rect 17099 28196 17133 28230
rect 17189 28196 17223 28230
rect 17279 28196 17313 28230
rect 17369 28196 17403 28230
rect 17459 28196 17493 28230
rect 16368 28112 16402 28146
rect 17555 28112 17589 28146
rect 16368 28022 16402 28056
rect 16368 27932 16402 27966
rect 16368 27842 16402 27876
rect 16368 27752 16402 27786
rect 16368 27662 16402 27696
rect 16368 27572 16402 27606
rect 16368 27482 16402 27516
rect 16368 27392 16402 27426
rect 16368 27302 16402 27336
rect 16368 27212 16402 27246
rect 16368 27122 16402 27156
rect 17555 28022 17589 28056
rect 17555 27932 17589 27966
rect 17555 27842 17589 27876
rect 17555 27752 17589 27786
rect 17555 27662 17589 27696
rect 17555 27572 17589 27606
rect 17555 27482 17589 27516
rect 17555 27392 17589 27426
rect 17555 27302 17589 27336
rect 17555 27212 17589 27246
rect 17555 27122 17589 27156
rect 16368 27032 16402 27066
rect 16469 27009 16503 27043
rect 16559 27009 16593 27043
rect 16649 27009 16683 27043
rect 16739 27009 16773 27043
rect 16829 27009 16863 27043
rect 16919 27009 16953 27043
rect 17009 27009 17043 27043
rect 17099 27009 17133 27043
rect 17189 27009 17223 27043
rect 17279 27009 17313 27043
rect 17369 27009 17403 27043
rect 17459 27009 17493 27043
rect 17555 27032 17589 27066
rect 13372 26825 13406 26963
rect 7552 26729 10352 26763
rect 10510 26729 13310 26763
rect 7456 26529 7490 26667
rect 10414 26529 10448 26667
rect 13372 26529 13406 26667
rect 7552 26433 10352 26467
rect 10510 26433 13310 26467
rect 7456 26233 7490 26371
rect 10414 26233 10448 26371
rect 13372 26233 13406 26371
rect 7552 26137 10352 26171
rect 10510 26137 13310 26171
rect 7456 25937 7490 26075
rect 10414 25937 10448 26075
rect 13372 25937 13406 26075
rect 7552 25841 10352 25875
rect 10510 25841 13310 25875
rect 7456 25641 7490 25779
rect 10414 25641 10448 25779
rect 13372 25641 13406 25779
rect 13781 26852 13815 26886
rect 13871 26852 13905 26886
rect 13961 26852 13995 26886
rect 14051 26852 14085 26886
rect 14141 26852 14175 26886
rect 14231 26852 14265 26886
rect 14321 26852 14355 26886
rect 14411 26852 14445 26886
rect 14501 26852 14535 26886
rect 14591 26852 14625 26886
rect 14681 26852 14715 26886
rect 14771 26852 14805 26886
rect 13680 26768 13714 26802
rect 14867 26768 14901 26802
rect 13680 26678 13714 26712
rect 13680 26588 13714 26622
rect 13680 26498 13714 26532
rect 13680 26408 13714 26442
rect 13680 26318 13714 26352
rect 13680 26228 13714 26262
rect 13680 26138 13714 26172
rect 13680 26048 13714 26082
rect 13680 25958 13714 25992
rect 13680 25868 13714 25902
rect 13680 25778 13714 25812
rect 14867 26678 14901 26712
rect 14867 26588 14901 26622
rect 14867 26498 14901 26532
rect 14867 26408 14901 26442
rect 14867 26318 14901 26352
rect 14867 26228 14901 26262
rect 14867 26138 14901 26172
rect 14867 26048 14901 26082
rect 14867 25958 14901 25992
rect 14867 25868 14901 25902
rect 14867 25778 14901 25812
rect 13680 25688 13714 25722
rect 13781 25665 13815 25699
rect 13871 25665 13905 25699
rect 13961 25665 13995 25699
rect 14051 25665 14085 25699
rect 14141 25665 14175 25699
rect 14231 25665 14265 25699
rect 14321 25665 14355 25699
rect 14411 25665 14445 25699
rect 14501 25665 14535 25699
rect 14591 25665 14625 25699
rect 14681 25665 14715 25699
rect 14771 25665 14805 25699
rect 14867 25688 14901 25722
rect 15125 26852 15159 26886
rect 15215 26852 15249 26886
rect 15305 26852 15339 26886
rect 15395 26852 15429 26886
rect 15485 26852 15519 26886
rect 15575 26852 15609 26886
rect 15665 26852 15699 26886
rect 15755 26852 15789 26886
rect 15845 26852 15879 26886
rect 15935 26852 15969 26886
rect 16025 26852 16059 26886
rect 16115 26852 16149 26886
rect 15024 26768 15058 26802
rect 16211 26768 16245 26802
rect 15024 26678 15058 26712
rect 15024 26588 15058 26622
rect 15024 26498 15058 26532
rect 15024 26408 15058 26442
rect 15024 26318 15058 26352
rect 15024 26228 15058 26262
rect 15024 26138 15058 26172
rect 15024 26048 15058 26082
rect 15024 25958 15058 25992
rect 15024 25868 15058 25902
rect 15024 25778 15058 25812
rect 16211 26678 16245 26712
rect 16211 26588 16245 26622
rect 16211 26498 16245 26532
rect 16211 26408 16245 26442
rect 16211 26318 16245 26352
rect 16211 26228 16245 26262
rect 16211 26138 16245 26172
rect 16211 26048 16245 26082
rect 16211 25958 16245 25992
rect 16211 25868 16245 25902
rect 16211 25778 16245 25812
rect 15024 25688 15058 25722
rect 15125 25665 15159 25699
rect 15215 25665 15249 25699
rect 15305 25665 15339 25699
rect 15395 25665 15429 25699
rect 15485 25665 15519 25699
rect 15575 25665 15609 25699
rect 15665 25665 15699 25699
rect 15755 25665 15789 25699
rect 15845 25665 15879 25699
rect 15935 25665 15969 25699
rect 16025 25665 16059 25699
rect 16115 25665 16149 25699
rect 16211 25688 16245 25722
rect 16469 26852 16503 26886
rect 16559 26852 16593 26886
rect 16649 26852 16683 26886
rect 16739 26852 16773 26886
rect 16829 26852 16863 26886
rect 16919 26852 16953 26886
rect 17009 26852 17043 26886
rect 17099 26852 17133 26886
rect 17189 26852 17223 26886
rect 17279 26852 17313 26886
rect 17369 26852 17403 26886
rect 17459 26852 17493 26886
rect 16368 26768 16402 26802
rect 17555 26768 17589 26802
rect 16368 26678 16402 26712
rect 16368 26588 16402 26622
rect 16368 26498 16402 26532
rect 16368 26408 16402 26442
rect 16368 26318 16402 26352
rect 16368 26228 16402 26262
rect 16368 26138 16402 26172
rect 16368 26048 16402 26082
rect 16368 25958 16402 25992
rect 16368 25868 16402 25902
rect 16368 25778 16402 25812
rect 17555 26678 17589 26712
rect 17555 26588 17589 26622
rect 17555 26498 17589 26532
rect 17555 26408 17589 26442
rect 17555 26318 17589 26352
rect 17555 26228 17589 26262
rect 17555 26138 17589 26172
rect 17555 26048 17589 26082
rect 17555 25958 17589 25992
rect 17555 25868 17589 25902
rect 17555 25778 17589 25812
rect 16368 25688 16402 25722
rect 16469 25665 16503 25699
rect 16559 25665 16593 25699
rect 16649 25665 16683 25699
rect 16739 25665 16773 25699
rect 16829 25665 16863 25699
rect 16919 25665 16953 25699
rect 17009 25665 17043 25699
rect 17099 25665 17133 25699
rect 17189 25665 17223 25699
rect 17279 25665 17313 25699
rect 17369 25665 17403 25699
rect 17459 25665 17493 25699
rect 17555 25688 17589 25722
rect 7552 25545 10352 25579
rect 10510 25545 13310 25579
rect 7456 25345 7490 25483
rect 10414 25345 10448 25483
rect 13372 25345 13406 25483
rect 7552 25249 10352 25283
rect 10510 25249 13310 25283
rect 7456 25049 7490 25187
rect 10414 25049 10448 25187
rect 13372 25049 13406 25187
rect 7552 24953 10352 24987
rect 10510 24953 13310 24987
rect 7456 24753 7490 24891
rect 10414 24753 10448 24891
rect 13372 24753 13406 24891
rect 7552 24657 10352 24691
rect 10510 24657 13310 24691
rect 13781 25508 13815 25542
rect 13871 25508 13905 25542
rect 13961 25508 13995 25542
rect 14051 25508 14085 25542
rect 14141 25508 14175 25542
rect 14231 25508 14265 25542
rect 14321 25508 14355 25542
rect 14411 25508 14445 25542
rect 14501 25508 14535 25542
rect 14591 25508 14625 25542
rect 14681 25508 14715 25542
rect 14771 25508 14805 25542
rect 13680 25424 13714 25458
rect 14867 25424 14901 25458
rect 13680 25334 13714 25368
rect 13680 25244 13714 25278
rect 13680 25154 13714 25188
rect 13680 25064 13714 25098
rect 13680 24974 13714 25008
rect 13680 24884 13714 24918
rect 13680 24794 13714 24828
rect 13680 24704 13714 24738
rect 13680 24614 13714 24648
rect 13680 24524 13714 24558
rect 13680 24434 13714 24468
rect 14867 25334 14901 25368
rect 14867 25244 14901 25278
rect 14867 25154 14901 25188
rect 14867 25064 14901 25098
rect 14867 24974 14901 25008
rect 14867 24884 14901 24918
rect 14867 24794 14901 24828
rect 14867 24704 14901 24738
rect 14867 24614 14901 24648
rect 14867 24524 14901 24558
rect 14867 24434 14901 24468
rect 13680 24344 13714 24378
rect 13781 24321 13815 24355
rect 13871 24321 13905 24355
rect 13961 24321 13995 24355
rect 14051 24321 14085 24355
rect 14141 24321 14175 24355
rect 14231 24321 14265 24355
rect 14321 24321 14355 24355
rect 14411 24321 14445 24355
rect 14501 24321 14535 24355
rect 14591 24321 14625 24355
rect 14681 24321 14715 24355
rect 14771 24321 14805 24355
rect 14867 24344 14901 24378
rect 15125 25508 15159 25542
rect 15215 25508 15249 25542
rect 15305 25508 15339 25542
rect 15395 25508 15429 25542
rect 15485 25508 15519 25542
rect 15575 25508 15609 25542
rect 15665 25508 15699 25542
rect 15755 25508 15789 25542
rect 15845 25508 15879 25542
rect 15935 25508 15969 25542
rect 16025 25508 16059 25542
rect 16115 25508 16149 25542
rect 15024 25424 15058 25458
rect 16211 25424 16245 25458
rect 15024 25334 15058 25368
rect 15024 25244 15058 25278
rect 15024 25154 15058 25188
rect 15024 25064 15058 25098
rect 15024 24974 15058 25008
rect 15024 24884 15058 24918
rect 15024 24794 15058 24828
rect 15024 24704 15058 24738
rect 15024 24614 15058 24648
rect 15024 24524 15058 24558
rect 15024 24434 15058 24468
rect 16211 25334 16245 25368
rect 16211 25244 16245 25278
rect 16211 25154 16245 25188
rect 16211 25064 16245 25098
rect 16211 24974 16245 25008
rect 16211 24884 16245 24918
rect 16211 24794 16245 24828
rect 16211 24704 16245 24738
rect 16211 24614 16245 24648
rect 16211 24524 16245 24558
rect 16211 24434 16245 24468
rect 15024 24344 15058 24378
rect 15125 24321 15159 24355
rect 15215 24321 15249 24355
rect 15305 24321 15339 24355
rect 15395 24321 15429 24355
rect 15485 24321 15519 24355
rect 15575 24321 15609 24355
rect 15665 24321 15699 24355
rect 15755 24321 15789 24355
rect 15845 24321 15879 24355
rect 15935 24321 15969 24355
rect 16025 24321 16059 24355
rect 16115 24321 16149 24355
rect 16211 24344 16245 24378
rect 16469 25508 16503 25542
rect 16559 25508 16593 25542
rect 16649 25508 16683 25542
rect 16739 25508 16773 25542
rect 16829 25508 16863 25542
rect 16919 25508 16953 25542
rect 17009 25508 17043 25542
rect 17099 25508 17133 25542
rect 17189 25508 17223 25542
rect 17279 25508 17313 25542
rect 17369 25508 17403 25542
rect 17459 25508 17493 25542
rect 16368 25424 16402 25458
rect 17555 25424 17589 25458
rect 16368 25334 16402 25368
rect 16368 25244 16402 25278
rect 16368 25154 16402 25188
rect 16368 25064 16402 25098
rect 16368 24974 16402 25008
rect 16368 24884 16402 24918
rect 16368 24794 16402 24828
rect 16368 24704 16402 24738
rect 16368 24614 16402 24648
rect 16368 24524 16402 24558
rect 16368 24434 16402 24468
rect 17555 25334 17589 25368
rect 17555 25244 17589 25278
rect 17555 25154 17589 25188
rect 17555 25064 17589 25098
rect 17555 24974 17589 25008
rect 17555 24884 17589 24918
rect 17555 24794 17589 24828
rect 17555 24704 17589 24738
rect 17555 24614 17589 24648
rect 17555 24524 17589 24558
rect 17555 24434 17589 24468
rect 16368 24344 16402 24378
rect 16469 24321 16503 24355
rect 16559 24321 16593 24355
rect 16649 24321 16683 24355
rect 16739 24321 16773 24355
rect 16829 24321 16863 24355
rect 16919 24321 16953 24355
rect 17009 24321 17043 24355
rect 17099 24321 17133 24355
rect 17189 24321 17223 24355
rect 17279 24321 17313 24355
rect 17369 24321 17403 24355
rect 17459 24321 17493 24355
rect 17555 24344 17589 24378
rect 14063 10793 14201 10827
rect 14359 10793 14497 10827
rect 14655 10793 14793 10827
rect 14951 10793 15089 10827
rect 15247 10793 15385 10827
rect 15543 10793 15681 10827
rect 15839 10793 15977 10827
rect 16135 10793 16273 10827
rect 13967 6731 14001 10731
rect 14263 6731 14297 10731
rect 14559 6731 14593 10731
rect 14855 6731 14889 10731
rect 15151 6731 15185 10731
rect 15447 6731 15481 10731
rect 15743 6731 15777 10731
rect 16039 6731 16073 10731
rect 16335 6731 16369 10731
rect 14063 6635 14201 6669
rect 14359 6635 14497 6669
rect 14655 6635 14793 6669
rect 14951 6635 15089 6669
rect 15247 6635 15385 6669
rect 15543 6635 15681 6669
rect 15839 6635 15977 6669
rect 16135 6635 16273 6669
rect 13967 2573 14001 6573
rect 14263 2573 14297 6573
rect 14559 2573 14593 6573
rect 14855 2573 14889 6573
rect 15151 2573 15185 6573
rect 15447 2573 15481 6573
rect 15743 2573 15777 6573
rect 16039 2573 16073 6573
rect 16335 2573 16369 6573
rect 18680 6335 18818 6369
rect 18976 6335 19114 6369
rect 19272 6335 19410 6369
rect 19568 6335 19706 6369
rect 14063 2477 14201 2511
rect 14359 2477 14497 2511
rect 14655 2477 14793 2511
rect 14951 2477 15089 2511
rect 15247 2477 15385 2511
rect 15543 2477 15681 2511
rect 15839 2477 15977 2511
rect 16135 2477 16273 2511
rect 18584 2573 18618 6273
rect 18880 2573 18914 6273
rect 19176 2573 19210 6273
rect 19472 2573 19506 6273
rect 19768 2573 19802 6273
rect 18680 2477 18818 2511
rect 18976 2477 19114 2511
rect 19272 2477 19410 2511
rect 19568 2477 19706 2511
<< nsubdiffcont >>
rect 13921 28046 13955 28080
rect 14011 28046 14045 28080
rect 14101 28046 14135 28080
rect 14191 28046 14225 28080
rect 14281 28046 14315 28080
rect 14371 28046 14405 28080
rect 14461 28046 14495 28080
rect 14551 28046 14585 28080
rect 14641 28046 14675 28080
rect 13829 27952 13863 27986
rect 13829 27862 13863 27896
rect 13829 27772 13863 27806
rect 13829 27682 13863 27716
rect 13829 27592 13863 27626
rect 13829 27502 13863 27536
rect 13829 27412 13863 27446
rect 13829 27322 13863 27356
rect 14719 27933 14753 27967
rect 14719 27843 14753 27877
rect 14719 27753 14753 27787
rect 14719 27663 14753 27697
rect 14719 27573 14753 27607
rect 14719 27483 14753 27517
rect 14719 27393 14753 27427
rect 14719 27303 14753 27337
rect 13829 27232 13863 27266
rect 14719 27213 14753 27247
rect 13887 27156 13921 27190
rect 13977 27156 14011 27190
rect 14067 27156 14101 27190
rect 14157 27156 14191 27190
rect 14247 27156 14281 27190
rect 14337 27156 14371 27190
rect 14427 27156 14461 27190
rect 14517 27156 14551 27190
rect 14607 27156 14641 27190
rect 15265 28046 15299 28080
rect 15355 28046 15389 28080
rect 15445 28046 15479 28080
rect 15535 28046 15569 28080
rect 15625 28046 15659 28080
rect 15715 28046 15749 28080
rect 15805 28046 15839 28080
rect 15895 28046 15929 28080
rect 15985 28046 16019 28080
rect 15173 27952 15207 27986
rect 15173 27862 15207 27896
rect 15173 27772 15207 27806
rect 15173 27682 15207 27716
rect 15173 27592 15207 27626
rect 15173 27502 15207 27536
rect 15173 27412 15207 27446
rect 15173 27322 15207 27356
rect 16063 27933 16097 27967
rect 16063 27843 16097 27877
rect 16063 27753 16097 27787
rect 16063 27663 16097 27697
rect 16063 27573 16097 27607
rect 16063 27483 16097 27517
rect 16063 27393 16097 27427
rect 16063 27303 16097 27337
rect 15173 27232 15207 27266
rect 16063 27213 16097 27247
rect 15231 27156 15265 27190
rect 15321 27156 15355 27190
rect 15411 27156 15445 27190
rect 15501 27156 15535 27190
rect 15591 27156 15625 27190
rect 15681 27156 15715 27190
rect 15771 27156 15805 27190
rect 15861 27156 15895 27190
rect 15951 27156 15985 27190
rect 16609 28046 16643 28080
rect 16699 28046 16733 28080
rect 16789 28046 16823 28080
rect 16879 28046 16913 28080
rect 16969 28046 17003 28080
rect 17059 28046 17093 28080
rect 17149 28046 17183 28080
rect 17239 28046 17273 28080
rect 17329 28046 17363 28080
rect 16517 27952 16551 27986
rect 16517 27862 16551 27896
rect 16517 27772 16551 27806
rect 16517 27682 16551 27716
rect 16517 27592 16551 27626
rect 16517 27502 16551 27536
rect 16517 27412 16551 27446
rect 16517 27322 16551 27356
rect 17407 27933 17441 27967
rect 17407 27843 17441 27877
rect 17407 27753 17441 27787
rect 17407 27663 17441 27697
rect 17407 27573 17441 27607
rect 17407 27483 17441 27517
rect 17407 27393 17441 27427
rect 17407 27303 17441 27337
rect 16517 27232 16551 27266
rect 17407 27213 17441 27247
rect 16575 27156 16609 27190
rect 16665 27156 16699 27190
rect 16755 27156 16789 27190
rect 16845 27156 16879 27190
rect 16935 27156 16969 27190
rect 17025 27156 17059 27190
rect 17115 27156 17149 27190
rect 17205 27156 17239 27190
rect 17295 27156 17329 27190
rect 13921 26702 13955 26736
rect 14011 26702 14045 26736
rect 14101 26702 14135 26736
rect 14191 26702 14225 26736
rect 14281 26702 14315 26736
rect 14371 26702 14405 26736
rect 14461 26702 14495 26736
rect 14551 26702 14585 26736
rect 14641 26702 14675 26736
rect 13829 26608 13863 26642
rect 13829 26518 13863 26552
rect 13829 26428 13863 26462
rect 13829 26338 13863 26372
rect 13829 26248 13863 26282
rect 13829 26158 13863 26192
rect 13829 26068 13863 26102
rect 13829 25978 13863 26012
rect 14719 26589 14753 26623
rect 14719 26499 14753 26533
rect 14719 26409 14753 26443
rect 14719 26319 14753 26353
rect 14719 26229 14753 26263
rect 14719 26139 14753 26173
rect 14719 26049 14753 26083
rect 14719 25959 14753 25993
rect 13829 25888 13863 25922
rect 14719 25869 14753 25903
rect 13887 25812 13921 25846
rect 13977 25812 14011 25846
rect 14067 25812 14101 25846
rect 14157 25812 14191 25846
rect 14247 25812 14281 25846
rect 14337 25812 14371 25846
rect 14427 25812 14461 25846
rect 14517 25812 14551 25846
rect 14607 25812 14641 25846
rect 15265 26702 15299 26736
rect 15355 26702 15389 26736
rect 15445 26702 15479 26736
rect 15535 26702 15569 26736
rect 15625 26702 15659 26736
rect 15715 26702 15749 26736
rect 15805 26702 15839 26736
rect 15895 26702 15929 26736
rect 15985 26702 16019 26736
rect 15173 26608 15207 26642
rect 15173 26518 15207 26552
rect 15173 26428 15207 26462
rect 15173 26338 15207 26372
rect 15173 26248 15207 26282
rect 15173 26158 15207 26192
rect 15173 26068 15207 26102
rect 15173 25978 15207 26012
rect 16063 26589 16097 26623
rect 16063 26499 16097 26533
rect 16063 26409 16097 26443
rect 16063 26319 16097 26353
rect 16063 26229 16097 26263
rect 16063 26139 16097 26173
rect 16063 26049 16097 26083
rect 16063 25959 16097 25993
rect 15173 25888 15207 25922
rect 16063 25869 16097 25903
rect 15231 25812 15265 25846
rect 15321 25812 15355 25846
rect 15411 25812 15445 25846
rect 15501 25812 15535 25846
rect 15591 25812 15625 25846
rect 15681 25812 15715 25846
rect 15771 25812 15805 25846
rect 15861 25812 15895 25846
rect 15951 25812 15985 25846
rect 16609 26702 16643 26736
rect 16699 26702 16733 26736
rect 16789 26702 16823 26736
rect 16879 26702 16913 26736
rect 16969 26702 17003 26736
rect 17059 26702 17093 26736
rect 17149 26702 17183 26736
rect 17239 26702 17273 26736
rect 17329 26702 17363 26736
rect 16517 26608 16551 26642
rect 16517 26518 16551 26552
rect 16517 26428 16551 26462
rect 16517 26338 16551 26372
rect 16517 26248 16551 26282
rect 16517 26158 16551 26192
rect 16517 26068 16551 26102
rect 16517 25978 16551 26012
rect 17407 26589 17441 26623
rect 17407 26499 17441 26533
rect 17407 26409 17441 26443
rect 17407 26319 17441 26353
rect 17407 26229 17441 26263
rect 17407 26139 17441 26173
rect 17407 26049 17441 26083
rect 17407 25959 17441 25993
rect 16517 25888 16551 25922
rect 17407 25869 17441 25903
rect 16575 25812 16609 25846
rect 16665 25812 16699 25846
rect 16755 25812 16789 25846
rect 16845 25812 16879 25846
rect 16935 25812 16969 25846
rect 17025 25812 17059 25846
rect 17115 25812 17149 25846
rect 17205 25812 17239 25846
rect 17295 25812 17329 25846
rect 13921 25358 13955 25392
rect 14011 25358 14045 25392
rect 14101 25358 14135 25392
rect 14191 25358 14225 25392
rect 14281 25358 14315 25392
rect 14371 25358 14405 25392
rect 14461 25358 14495 25392
rect 14551 25358 14585 25392
rect 14641 25358 14675 25392
rect 13829 25264 13863 25298
rect 13829 25174 13863 25208
rect 13829 25084 13863 25118
rect 13829 24994 13863 25028
rect 13829 24904 13863 24938
rect 13829 24814 13863 24848
rect 13829 24724 13863 24758
rect 13829 24634 13863 24668
rect 14719 25245 14753 25279
rect 14719 25155 14753 25189
rect 14719 25065 14753 25099
rect 14719 24975 14753 25009
rect 14719 24885 14753 24919
rect 14719 24795 14753 24829
rect 14719 24705 14753 24739
rect 14719 24615 14753 24649
rect 13829 24544 13863 24578
rect 14719 24525 14753 24559
rect 13887 24468 13921 24502
rect 13977 24468 14011 24502
rect 14067 24468 14101 24502
rect 14157 24468 14191 24502
rect 14247 24468 14281 24502
rect 14337 24468 14371 24502
rect 14427 24468 14461 24502
rect 14517 24468 14551 24502
rect 14607 24468 14641 24502
rect 15265 25358 15299 25392
rect 15355 25358 15389 25392
rect 15445 25358 15479 25392
rect 15535 25358 15569 25392
rect 15625 25358 15659 25392
rect 15715 25358 15749 25392
rect 15805 25358 15839 25392
rect 15895 25358 15929 25392
rect 15985 25358 16019 25392
rect 15173 25264 15207 25298
rect 15173 25174 15207 25208
rect 15173 25084 15207 25118
rect 15173 24994 15207 25028
rect 15173 24904 15207 24938
rect 15173 24814 15207 24848
rect 15173 24724 15207 24758
rect 15173 24634 15207 24668
rect 16063 25245 16097 25279
rect 16063 25155 16097 25189
rect 16063 25065 16097 25099
rect 16063 24975 16097 25009
rect 16063 24885 16097 24919
rect 16063 24795 16097 24829
rect 16063 24705 16097 24739
rect 16063 24615 16097 24649
rect 15173 24544 15207 24578
rect 16063 24525 16097 24559
rect 15231 24468 15265 24502
rect 15321 24468 15355 24502
rect 15411 24468 15445 24502
rect 15501 24468 15535 24502
rect 15591 24468 15625 24502
rect 15681 24468 15715 24502
rect 15771 24468 15805 24502
rect 15861 24468 15895 24502
rect 15951 24468 15985 24502
rect 16609 25358 16643 25392
rect 16699 25358 16733 25392
rect 16789 25358 16823 25392
rect 16879 25358 16913 25392
rect 16969 25358 17003 25392
rect 17059 25358 17093 25392
rect 17149 25358 17183 25392
rect 17239 25358 17273 25392
rect 17329 25358 17363 25392
rect 16517 25264 16551 25298
rect 16517 25174 16551 25208
rect 16517 25084 16551 25118
rect 16517 24994 16551 25028
rect 16517 24904 16551 24938
rect 16517 24814 16551 24848
rect 16517 24724 16551 24758
rect 16517 24634 16551 24668
rect 17407 25245 17441 25279
rect 17407 25155 17441 25189
rect 17407 25065 17441 25099
rect 17407 24975 17441 25009
rect 17407 24885 17441 24919
rect 17407 24795 17441 24829
rect 17407 24705 17441 24739
rect 17407 24615 17441 24649
rect 16517 24544 16551 24578
rect 17407 24525 17441 24559
rect 16575 24468 16609 24502
rect 16665 24468 16699 24502
rect 16755 24468 16789 24502
rect 16845 24468 16879 24502
rect 16935 24468 16969 24502
rect 17025 24468 17059 24502
rect 17115 24468 17149 24502
rect 17205 24468 17239 24502
rect 17295 24468 17329 24502
<< mvpsubdiffcont >>
rect 6038 24202 6366 24236
rect 6524 24202 6852 24236
rect 7010 24202 7338 24236
rect 7496 24202 7824 24236
rect 7982 24202 8310 24236
rect 8468 24202 8796 24236
rect 8954 24202 9282 24236
rect 9440 24202 9768 24236
rect 9926 24202 10254 24236
rect 10412 24202 10740 24236
rect 5942 19972 5976 24140
rect 6428 19972 6462 24140
rect 6914 19972 6948 24140
rect 7400 19972 7434 24140
rect 7886 19972 7920 24140
rect 8372 19972 8406 24140
rect 8858 19972 8892 24140
rect 9344 19972 9378 24140
rect 9830 19972 9864 24140
rect 10316 19972 10350 24140
rect 10802 19972 10836 24140
rect 15759 23795 19927 23829
rect 11303 23395 15471 23429
rect 11207 22505 11241 23333
rect 15533 22505 15567 23333
rect 11303 22409 15471 22443
rect 15663 22505 15697 23733
rect 19989 22505 20023 23733
rect 15759 22409 19927 22443
rect 11310 22123 15478 22157
rect 11214 20833 11248 22061
rect 15540 20833 15574 22061
rect 15759 22123 19927 22157
rect 15663 21233 15697 22061
rect 19989 21233 20023 22061
rect 15759 21137 19927 21171
rect 11310 20737 15478 20771
rect 6038 19876 6366 19910
rect 6524 19876 6852 19910
rect 7010 19876 7338 19910
rect 7496 19876 7824 19910
rect 7982 19876 8310 19910
rect 8468 19876 8796 19910
rect 8954 19876 9282 19910
rect 9440 19876 9768 19910
rect 9926 19876 10254 19910
rect 10412 19876 10740 19910
rect 11379 9826 11647 9860
rect 11283 9336 11317 9764
rect 11709 9336 11743 9764
rect 11379 9240 11647 9274
rect 11935 9826 12203 9860
rect 11839 9336 11873 9764
rect 12265 9336 12299 9764
rect 11935 9240 12203 9274
rect 12491 9826 12759 9860
rect 12395 9336 12429 9764
rect 12821 9336 12855 9764
rect 12491 9240 12759 9274
rect 13047 9826 13315 9860
rect 12951 9336 12985 9764
rect 13377 9336 13411 9764
rect 13047 9240 13315 9274
rect 5427 8575 6795 8609
rect 5331 8085 5365 8513
rect 6857 8085 6891 8513
rect 5427 7989 6795 8023
rect 7083 8575 8451 8609
rect 6987 8085 7021 8513
rect 8513 8085 8547 8513
rect 7083 7989 8451 8023
rect 9013 8575 9621 8609
rect 8917 8085 8951 8513
rect 9683 8085 9717 8513
rect 9013 7989 9621 8023
rect 9985 8576 10593 8610
rect 9889 8086 9923 8514
rect 10655 8086 10689 8514
rect 9985 7990 10593 8024
rect 5427 7859 6795 7893
rect 5331 7369 5365 7797
rect 6857 7369 6891 7797
rect 5427 7273 6795 7307
rect 7083 7859 8451 7893
rect 6987 7369 7021 7797
rect 8513 7369 8547 7797
rect 7083 7273 8451 7307
rect 5427 7143 6795 7177
rect 5331 6653 5365 7081
rect 6857 6653 6891 7081
rect 5427 6557 6795 6591
rect 7083 7143 8451 7177
rect 6987 6653 7021 7081
rect 8513 6653 8547 7081
rect 7083 6557 8451 6591
rect 16571 9864 20157 9898
rect 16475 7574 16509 9802
rect 20219 7574 20253 9802
rect 16571 7478 20157 7512
rect 21623 8045 23851 8079
rect 5427 6427 6795 6461
rect 5331 5937 5365 6365
rect 6857 5937 6891 6365
rect 5427 5841 6795 5875
rect 7083 6427 8451 6461
rect 6987 5937 7021 6365
rect 8513 5937 8547 6365
rect 7083 5841 8451 5875
rect 16567 7277 16995 7311
rect 17153 7277 17581 7311
rect 17739 7277 18167 7311
rect 16471 5047 16505 7215
rect 17057 5047 17091 7215
rect 17643 5047 17677 7215
rect 18229 5047 18263 7215
rect 16567 4951 16995 4985
rect 17153 4951 17581 4985
rect 17739 4951 18167 4985
rect 16567 4815 16995 4849
rect 17153 4815 17581 4849
rect 17739 4815 18167 4849
rect 16471 2585 16505 4753
rect 17057 2585 17091 4753
rect 17643 2585 17677 4753
rect 18229 2585 18263 4753
rect 16567 2489 16995 2523
rect 17153 2489 17581 2523
rect 17739 2489 18167 2523
rect 21527 6015 21561 7983
rect 23913 6015 23947 7983
rect 21623 5919 23851 5953
rect 21623 5795 23851 5829
rect 21527 3765 21561 5733
rect 23913 3765 23947 5733
rect 21623 3669 23851 3703
rect 24552 3937 26780 3971
rect 21408 3103 24098 3137
rect 21312 1813 21346 3041
rect 24160 1813 24194 3041
rect 24456 1907 24490 3875
rect 26842 1907 26876 3875
rect 24552 1811 26780 1845
rect 21408 1717 24098 1751
<< mvnsubdiffcont >>
rect 6195 31103 8363 31137
rect 8521 31103 10689 31137
rect 6099 30595 6133 31041
rect 8425 30595 8459 31041
rect 10751 30595 10785 31041
rect 6195 30499 8363 30533
rect 8521 30499 10689 30533
rect 6320 19236 10488 19270
rect 6224 18092 6258 19174
rect 10550 18092 10584 19174
rect 6320 17996 10488 18030
rect 11408 19236 15576 19270
rect 15734 19236 19902 19270
rect 6320 17836 10488 17870
rect 6224 16928 6258 17774
rect 10550 16928 10584 17774
rect 6320 16832 10488 16866
rect 11312 16928 11346 19174
rect 15638 16928 15672 19174
rect 19964 16928 19998 19174
rect 11408 16832 15576 16866
rect 15734 16832 19902 16866
rect 8330 15032 10488 15066
rect 8234 14524 8268 14970
rect 10550 14524 10584 14970
rect 8330 14428 10488 14462
rect 11312 14524 11346 16770
rect 15638 14524 15672 16770
rect 19964 14524 19998 16770
rect 20776 18868 21122 18902
rect 21280 18868 21626 18902
rect 20680 14638 20714 18806
rect 21184 14638 21218 18806
rect 21688 14638 21722 18806
rect 20776 14542 21122 14576
rect 21280 14542 21626 14576
rect 11408 14428 15576 14462
rect 15734 14428 19902 14462
rect 8035 12508 10213 12542
rect 7939 12000 7973 12446
rect 10275 12000 10309 12446
rect 8035 11904 10213 11938
rect 6035 11745 10203 11779
rect 5939 11037 5973 11683
rect 10265 11037 10299 11683
rect 6035 10941 10203 10975
rect 11973 11015 12757 11049
rect 6147 10759 6795 10793
rect 6051 9951 6085 10697
rect 6857 9951 6891 10697
rect 6147 9855 6795 9889
rect 7083 10759 7731 10793
rect 6987 9951 7021 10697
rect 7793 9951 7827 10697
rect 7083 9855 7731 9889
rect 9013 10777 9661 10811
rect 8917 9969 8951 10715
rect 9723 9969 9757 10715
rect 9013 9873 9661 9907
rect 9945 10777 10593 10811
rect 9849 9969 9883 10715
rect 10655 9969 10689 10715
rect 11913 10533 11947 10989
rect 12783 10533 12817 10989
rect 11973 10473 12757 10507
rect 9945 9873 10593 9907
rect 6147 9717 6795 9751
rect 6051 8909 6085 9655
rect 6857 8909 6891 9655
rect 6147 8813 6795 8847
rect 7083 9717 7731 9751
rect 6987 8909 7021 9655
rect 7793 8909 7827 9655
rect 7083 8813 7731 8847
rect 9013 9692 9661 9726
rect 8917 8884 8951 9630
rect 9723 8884 9757 9630
rect 9013 8788 9661 8822
rect 9945 9692 10593 9726
rect 9849 8884 9883 9630
rect 10655 8884 10689 9630
rect 9945 8788 10593 8822
rect 24708 8045 25754 8079
rect 24612 7615 24646 7983
rect 25816 7615 25850 7983
rect 24708 7519 25754 7553
rect 24708 7339 26654 7373
rect 24612 5103 24646 7277
rect 26716 5103 26750 7277
rect 24708 5007 26654 5041
<< poly >>
rect 6279 30999 8279 31015
rect 6279 30965 6295 30999
rect 8263 30965 8279 30999
rect 6279 30918 8279 30965
rect 6279 30671 8279 30718
rect 6279 30637 6295 30671
rect 8263 30637 8279 30671
rect 6279 30621 8279 30637
rect 8605 30999 10605 31015
rect 8605 30965 8621 30999
rect 10589 30965 10605 30999
rect 8605 30918 10605 30965
rect 8605 30671 10605 30718
rect 8605 30637 8621 30671
rect 10589 30637 10605 30671
rect 8605 30621 10605 30637
rect 6064 24040 6152 24056
rect 6064 20072 6080 24040
rect 6114 20072 6152 24040
rect 6064 20056 6152 20072
rect 6252 24040 6340 24056
rect 6252 20072 6290 24040
rect 6324 20072 6340 24040
rect 6252 20056 6340 20072
rect 6550 24040 6638 24056
rect 6550 20072 6566 24040
rect 6600 20072 6638 24040
rect 6550 20056 6638 20072
rect 6738 24040 6826 24056
rect 6738 20072 6776 24040
rect 6810 20072 6826 24040
rect 6738 20056 6826 20072
rect 7036 24040 7124 24056
rect 7036 20072 7052 24040
rect 7086 20072 7124 24040
rect 7036 20056 7124 20072
rect 7224 24040 7312 24056
rect 7224 20072 7262 24040
rect 7296 20072 7312 24040
rect 7224 20056 7312 20072
rect 7522 24040 7610 24056
rect 7522 20072 7538 24040
rect 7572 20072 7610 24040
rect 7522 20056 7610 20072
rect 7710 24040 7798 24056
rect 7710 20072 7748 24040
rect 7782 20072 7798 24040
rect 7710 20056 7798 20072
rect 8008 24040 8096 24056
rect 8008 20072 8024 24040
rect 8058 20072 8096 24040
rect 8008 20056 8096 20072
rect 8196 24040 8284 24056
rect 8196 20072 8234 24040
rect 8268 20072 8284 24040
rect 8196 20056 8284 20072
rect 8494 24040 8582 24056
rect 8494 20072 8510 24040
rect 8544 20072 8582 24040
rect 8494 20056 8582 20072
rect 8682 24040 8770 24056
rect 8682 20072 8720 24040
rect 8754 20072 8770 24040
rect 8682 20056 8770 20072
rect 8980 24040 9068 24056
rect 8980 20072 8996 24040
rect 9030 20072 9068 24040
rect 8980 20056 9068 20072
rect 9168 24040 9256 24056
rect 9168 20072 9206 24040
rect 9240 20072 9256 24040
rect 9168 20056 9256 20072
rect 9466 24040 9554 24056
rect 9466 20072 9482 24040
rect 9516 20072 9554 24040
rect 9466 20056 9554 20072
rect 9654 24040 9742 24056
rect 9654 20072 9692 24040
rect 9726 20072 9742 24040
rect 9654 20056 9742 20072
rect 9952 24040 10040 24056
rect 9952 20072 9968 24040
rect 10002 20072 10040 24040
rect 9952 20056 10040 20072
rect 10140 24040 10228 24056
rect 10140 20072 10178 24040
rect 10212 20072 10228 24040
rect 10140 20056 10228 20072
rect 10438 24040 10526 24056
rect 10438 20072 10454 24040
rect 10488 20072 10526 24040
rect 10438 20056 10526 20072
rect 10626 24040 10714 24056
rect 10626 20072 10664 24040
rect 10698 20072 10714 24040
rect 10626 20056 10714 20072
rect 11387 23291 15387 23307
rect 11387 23257 11403 23291
rect 15371 23257 15387 23291
rect 11387 23219 15387 23257
rect 11387 22581 15387 22619
rect 11387 22547 11403 22581
rect 15371 22547 15387 22581
rect 11387 22531 15387 22547
rect 15843 23691 19843 23707
rect 15843 23657 15859 23691
rect 19827 23657 19843 23691
rect 15843 23619 19843 23657
rect 15843 22581 19843 22619
rect 15843 22547 15859 22581
rect 19827 22547 19843 22581
rect 15843 22531 19843 22547
rect 11394 22019 15394 22035
rect 11394 21985 11410 22019
rect 15378 21985 15394 22019
rect 11394 21947 15394 21985
rect 11394 20909 15394 20947
rect 11394 20875 11410 20909
rect 15378 20875 15394 20909
rect 11394 20859 15394 20875
rect 15843 22019 19843 22035
rect 15843 21985 15859 22019
rect 19827 21985 19843 22019
rect 15843 21947 19843 21985
rect 15843 21309 19843 21347
rect 15843 21275 15859 21309
rect 19827 21275 19843 21309
rect 15843 21259 19843 21275
rect 6404 19132 10404 19148
rect 6404 19098 6420 19132
rect 10388 19098 10404 19132
rect 6404 19051 10404 19098
rect 6404 18704 10404 18751
rect 6404 18670 6420 18704
rect 10388 18670 10404 18704
rect 6404 18654 10404 18670
rect 6404 18596 10404 18612
rect 6404 18562 6420 18596
rect 10388 18562 10404 18596
rect 6404 18515 10404 18562
rect 6404 18168 10404 18215
rect 6404 18134 6420 18168
rect 10388 18134 10404 18168
rect 6404 18118 10404 18134
rect 6404 17732 10404 17748
rect 6404 17698 6420 17732
rect 10388 17698 10404 17732
rect 6404 17651 10404 17698
rect 6404 17004 10404 17051
rect 6404 16970 6420 17004
rect 10388 16970 10404 17004
rect 6404 16954 10404 16970
rect 11492 19132 15492 19148
rect 11492 19098 11508 19132
rect 15476 19098 15492 19132
rect 11492 19051 15492 19098
rect 11492 17004 15492 17051
rect 11492 16970 11508 17004
rect 15476 16970 15492 17004
rect 11492 16954 15492 16970
rect 15818 19132 19818 19148
rect 15818 19098 15834 19132
rect 19802 19098 19818 19132
rect 15818 19051 19818 19098
rect 15818 17004 19818 17051
rect 15818 16970 15834 17004
rect 19802 16970 19818 17004
rect 15818 16954 19818 16970
rect 8414 14928 10404 14944
rect 8414 14894 8430 14928
rect 10388 14894 10404 14928
rect 8414 14847 10404 14894
rect 8414 14600 10404 14647
rect 8414 14566 8430 14600
rect 10388 14566 10404 14600
rect 8414 14550 10404 14566
rect 11492 16728 15492 16744
rect 11492 16694 11508 16728
rect 15476 16694 15492 16728
rect 11492 16647 15492 16694
rect 11492 14600 15492 14647
rect 11492 14566 11508 14600
rect 15476 14566 15492 14600
rect 11492 14550 15492 14566
rect 15818 16728 19818 16744
rect 15818 16694 15834 16728
rect 19802 16694 19818 16728
rect 15818 16647 19818 16694
rect 15818 14600 19818 14647
rect 15818 14566 15834 14600
rect 19802 14566 19818 14600
rect 15818 14550 19818 14566
rect 20802 18706 20899 18722
rect 20802 14738 20818 18706
rect 20852 14738 20899 18706
rect 20802 14722 20899 14738
rect 20999 18706 21096 18722
rect 20999 14738 21046 18706
rect 21080 14738 21096 18706
rect 20999 14722 21096 14738
rect 21306 18706 21403 18722
rect 21306 14738 21322 18706
rect 21356 14738 21403 18706
rect 21306 14722 21403 14738
rect 21503 18706 21600 18722
rect 21503 14738 21550 18706
rect 21584 14738 21600 18706
rect 21503 14722 21600 14738
rect 8119 12404 10129 12420
rect 8119 12370 8135 12404
rect 10113 12370 10129 12404
rect 8119 12323 10129 12370
rect 8119 12076 10129 12123
rect 8119 12042 8135 12076
rect 10113 12042 10129 12076
rect 8119 12026 10129 12042
rect 6119 11641 10119 11657
rect 6119 11607 6135 11641
rect 10103 11607 10119 11641
rect 6119 11560 10119 11607
rect 6119 11113 10119 11160
rect 6119 11079 6135 11113
rect 10103 11079 10119 11113
rect 6119 11063 10119 11079
rect 6231 10655 6711 10671
rect 6231 10621 6247 10655
rect 6695 10621 6711 10655
rect 6231 10574 6711 10621
rect 6231 10027 6711 10074
rect 6231 9993 6247 10027
rect 6695 9993 6711 10027
rect 6231 9977 6711 9993
rect 7167 10655 7647 10671
rect 7167 10621 7183 10655
rect 7631 10621 7647 10655
rect 7167 10574 7647 10621
rect 7167 10027 7647 10074
rect 7167 9993 7183 10027
rect 7631 9993 7647 10027
rect 7167 9977 7647 9993
rect 9097 10673 9577 10689
rect 9097 10639 9113 10673
rect 9561 10639 9577 10673
rect 9097 10592 9577 10639
rect 9097 10045 9577 10092
rect 9097 10011 9113 10045
rect 9561 10011 9577 10045
rect 9097 9995 9577 10011
rect 10029 10673 10509 10689
rect 10029 10639 10045 10673
rect 10493 10639 10509 10673
rect 10029 10592 10509 10639
rect 10029 10045 10509 10092
rect 10029 10011 10045 10045
rect 10493 10011 10509 10045
rect 10029 9995 10509 10011
rect 12079 10946 12179 10962
rect 12079 10912 12095 10946
rect 12163 10912 12179 10946
rect 12079 10865 12179 10912
rect 12237 10946 12337 10962
rect 12237 10912 12253 10946
rect 12321 10912 12337 10946
rect 12237 10865 12337 10912
rect 12395 10946 12495 10962
rect 12395 10912 12411 10946
rect 12479 10912 12495 10946
rect 12395 10865 12495 10912
rect 12553 10946 12653 10962
rect 12553 10912 12569 10946
rect 12637 10912 12653 10946
rect 12553 10865 12653 10912
rect 12079 10618 12179 10665
rect 12079 10584 12095 10618
rect 12163 10584 12179 10618
rect 12079 10568 12179 10584
rect 12237 10618 12337 10665
rect 12237 10584 12253 10618
rect 12321 10584 12337 10618
rect 12237 10568 12337 10584
rect 12395 10618 12495 10665
rect 12395 10584 12411 10618
rect 12479 10584 12495 10618
rect 12395 10568 12495 10584
rect 12553 10618 12653 10665
rect 12553 10584 12569 10618
rect 12637 10584 12653 10618
rect 12553 10568 12653 10584
rect 6231 9613 6711 9629
rect 6231 9579 6247 9613
rect 6695 9579 6711 9613
rect 6231 9532 6711 9579
rect 6231 8985 6711 9032
rect 6231 8951 6247 8985
rect 6695 8951 6711 8985
rect 6231 8935 6711 8951
rect 7167 9613 7647 9629
rect 7167 9579 7183 9613
rect 7631 9579 7647 9613
rect 7167 9532 7647 9579
rect 7167 8985 7647 9032
rect 7167 8951 7183 8985
rect 7631 8951 7647 8985
rect 7167 8935 7647 8951
rect 9097 9588 9577 9604
rect 9097 9554 9113 9588
rect 9561 9554 9577 9588
rect 9097 9507 9577 9554
rect 9097 8960 9577 9007
rect 9097 8926 9113 8960
rect 9561 8926 9577 8960
rect 9097 8910 9577 8926
rect 10029 9588 10509 9604
rect 10029 9554 10045 9588
rect 10493 9554 10509 9588
rect 10029 9507 10509 9554
rect 10029 8960 10509 9007
rect 10029 8926 10045 8960
rect 10493 8926 10509 8960
rect 10029 8910 10509 8926
rect 11463 9722 11563 9738
rect 11463 9688 11479 9722
rect 11547 9688 11563 9722
rect 11463 9650 11563 9688
rect 11463 9412 11563 9450
rect 11463 9378 11479 9412
rect 11547 9378 11563 9412
rect 11463 9362 11563 9378
rect 12019 9722 12119 9738
rect 12019 9688 12035 9722
rect 12103 9688 12119 9722
rect 12019 9650 12119 9688
rect 12019 9412 12119 9450
rect 12019 9378 12035 9412
rect 12103 9378 12119 9412
rect 12019 9362 12119 9378
rect 12575 9722 12675 9738
rect 12575 9688 12591 9722
rect 12659 9688 12675 9722
rect 12575 9650 12675 9688
rect 12575 9412 12675 9450
rect 12575 9378 12591 9412
rect 12659 9378 12675 9412
rect 12575 9362 12675 9378
rect 13131 9722 13231 9738
rect 13131 9688 13147 9722
rect 13215 9688 13231 9722
rect 13131 9650 13231 9688
rect 13131 9412 13231 9450
rect 13131 9378 13147 9412
rect 13215 9378 13231 9412
rect 13131 9362 13231 9378
rect 5511 8471 6711 8487
rect 5511 8437 5527 8471
rect 6695 8437 6711 8471
rect 5511 8399 6711 8437
rect 5511 8161 6711 8199
rect 5511 8127 5527 8161
rect 6695 8127 6711 8161
rect 5511 8111 6711 8127
rect 7167 8471 8367 8487
rect 7167 8437 7183 8471
rect 8351 8437 8367 8471
rect 7167 8399 8367 8437
rect 7167 8161 8367 8199
rect 7167 8127 7183 8161
rect 8351 8127 8367 8161
rect 7167 8111 8367 8127
rect 9097 8471 9537 8487
rect 9097 8437 9113 8471
rect 9521 8437 9537 8471
rect 9097 8399 9537 8437
rect 9097 8161 9537 8199
rect 9097 8127 9113 8161
rect 9521 8127 9537 8161
rect 9097 8111 9537 8127
rect 10069 8472 10509 8488
rect 10069 8438 10085 8472
rect 10493 8438 10509 8472
rect 10069 8400 10509 8438
rect 10069 8162 10509 8200
rect 10069 8128 10085 8162
rect 10493 8128 10509 8162
rect 10069 8112 10509 8128
rect 5511 7755 6711 7771
rect 5511 7721 5527 7755
rect 6695 7721 6711 7755
rect 5511 7683 6711 7721
rect 5511 7445 6711 7483
rect 5511 7411 5527 7445
rect 6695 7411 6711 7445
rect 5511 7395 6711 7411
rect 7167 7755 8367 7771
rect 7167 7721 7183 7755
rect 8351 7721 8367 7755
rect 7167 7683 8367 7721
rect 7167 7445 8367 7483
rect 7167 7411 7183 7445
rect 8351 7411 8367 7445
rect 7167 7395 8367 7411
rect 5511 7039 6711 7055
rect 5511 7005 5527 7039
rect 6695 7005 6711 7039
rect 5511 6967 6711 7005
rect 5511 6729 6711 6767
rect 5511 6695 5527 6729
rect 6695 6695 6711 6729
rect 5511 6679 6711 6695
rect 7167 7039 8367 7055
rect 7167 7005 7183 7039
rect 8351 7005 8367 7039
rect 7167 6967 8367 7005
rect 7167 6729 8367 6767
rect 7167 6695 7183 6729
rect 8351 6695 8367 6729
rect 7167 6679 8367 6695
rect 16655 9760 16755 9776
rect 16655 9726 16671 9760
rect 16739 9726 16755 9760
rect 16655 9688 16755 9726
rect 16813 9760 16913 9776
rect 16813 9726 16829 9760
rect 16897 9726 16913 9760
rect 16813 9688 16913 9726
rect 16971 9760 17071 9776
rect 16971 9726 16987 9760
rect 17055 9726 17071 9760
rect 16971 9688 17071 9726
rect 17129 9760 17229 9776
rect 17129 9726 17145 9760
rect 17213 9726 17229 9760
rect 17129 9688 17229 9726
rect 17287 9760 17387 9776
rect 17287 9726 17303 9760
rect 17371 9726 17387 9760
rect 17287 9688 17387 9726
rect 17445 9760 17545 9776
rect 17445 9726 17461 9760
rect 17529 9726 17545 9760
rect 17445 9688 17545 9726
rect 17603 9760 17703 9776
rect 17603 9726 17619 9760
rect 17687 9726 17703 9760
rect 17603 9688 17703 9726
rect 17761 9760 17861 9776
rect 17761 9726 17777 9760
rect 17845 9726 17861 9760
rect 17761 9688 17861 9726
rect 17919 9760 18019 9776
rect 17919 9726 17935 9760
rect 18003 9726 18019 9760
rect 17919 9688 18019 9726
rect 18077 9760 18177 9776
rect 18077 9726 18093 9760
rect 18161 9726 18177 9760
rect 18077 9688 18177 9726
rect 18235 9760 18335 9776
rect 18235 9726 18251 9760
rect 18319 9726 18335 9760
rect 18235 9688 18335 9726
rect 18393 9760 18493 9776
rect 18393 9726 18409 9760
rect 18477 9726 18493 9760
rect 18393 9688 18493 9726
rect 18551 9760 18651 9776
rect 18551 9726 18567 9760
rect 18635 9726 18651 9760
rect 18551 9688 18651 9726
rect 18709 9760 18809 9776
rect 18709 9726 18725 9760
rect 18793 9726 18809 9760
rect 18709 9688 18809 9726
rect 18867 9760 18967 9776
rect 18867 9726 18883 9760
rect 18951 9726 18967 9760
rect 18867 9688 18967 9726
rect 19025 9760 19125 9776
rect 19025 9726 19041 9760
rect 19109 9726 19125 9760
rect 19025 9688 19125 9726
rect 19183 9760 19283 9776
rect 19183 9726 19199 9760
rect 19267 9726 19283 9760
rect 19183 9688 19283 9726
rect 19341 9760 19441 9776
rect 19341 9726 19357 9760
rect 19425 9726 19441 9760
rect 19341 9688 19441 9726
rect 19499 9760 19599 9776
rect 19499 9726 19515 9760
rect 19583 9726 19599 9760
rect 19499 9688 19599 9726
rect 19657 9760 19757 9776
rect 19657 9726 19673 9760
rect 19741 9726 19757 9760
rect 19657 9688 19757 9726
rect 19815 9760 19915 9776
rect 19815 9726 19831 9760
rect 19899 9726 19915 9760
rect 19815 9688 19915 9726
rect 19973 9760 20073 9776
rect 19973 9726 19989 9760
rect 20057 9726 20073 9760
rect 19973 9688 20073 9726
rect 16655 7650 16755 7688
rect 16655 7616 16671 7650
rect 16739 7616 16755 7650
rect 16655 7600 16755 7616
rect 16813 7650 16913 7688
rect 16813 7616 16829 7650
rect 16897 7616 16913 7650
rect 16813 7600 16913 7616
rect 16971 7650 17071 7688
rect 16971 7616 16987 7650
rect 17055 7616 17071 7650
rect 16971 7600 17071 7616
rect 17129 7650 17229 7688
rect 17129 7616 17145 7650
rect 17213 7616 17229 7650
rect 17129 7600 17229 7616
rect 17287 7650 17387 7688
rect 17287 7616 17303 7650
rect 17371 7616 17387 7650
rect 17287 7600 17387 7616
rect 17445 7650 17545 7688
rect 17445 7616 17461 7650
rect 17529 7616 17545 7650
rect 17445 7600 17545 7616
rect 17603 7650 17703 7688
rect 17603 7616 17619 7650
rect 17687 7616 17703 7650
rect 17603 7600 17703 7616
rect 17761 7650 17861 7688
rect 17761 7616 17777 7650
rect 17845 7616 17861 7650
rect 17761 7600 17861 7616
rect 17919 7650 18019 7688
rect 17919 7616 17935 7650
rect 18003 7616 18019 7650
rect 17919 7600 18019 7616
rect 18077 7650 18177 7688
rect 18077 7616 18093 7650
rect 18161 7616 18177 7650
rect 18077 7600 18177 7616
rect 18235 7650 18335 7688
rect 18235 7616 18251 7650
rect 18319 7616 18335 7650
rect 18235 7600 18335 7616
rect 18393 7650 18493 7688
rect 18393 7616 18409 7650
rect 18477 7616 18493 7650
rect 18393 7600 18493 7616
rect 18551 7650 18651 7688
rect 18551 7616 18567 7650
rect 18635 7616 18651 7650
rect 18551 7600 18651 7616
rect 18709 7650 18809 7688
rect 18709 7616 18725 7650
rect 18793 7616 18809 7650
rect 18709 7600 18809 7616
rect 18867 7650 18967 7688
rect 18867 7616 18883 7650
rect 18951 7616 18967 7650
rect 18867 7600 18967 7616
rect 19025 7650 19125 7688
rect 19025 7616 19041 7650
rect 19109 7616 19125 7650
rect 19025 7600 19125 7616
rect 19183 7650 19283 7688
rect 19183 7616 19199 7650
rect 19267 7616 19283 7650
rect 19183 7600 19283 7616
rect 19341 7650 19441 7688
rect 19341 7616 19357 7650
rect 19425 7616 19441 7650
rect 19341 7600 19441 7616
rect 19499 7650 19599 7688
rect 19499 7616 19515 7650
rect 19583 7616 19599 7650
rect 19499 7600 19599 7616
rect 19657 7650 19757 7688
rect 19657 7616 19673 7650
rect 19741 7616 19757 7650
rect 19657 7600 19757 7616
rect 19815 7650 19915 7688
rect 19815 7616 19831 7650
rect 19899 7616 19915 7650
rect 19815 7600 19915 7616
rect 19973 7650 20073 7688
rect 19973 7616 19989 7650
rect 20057 7616 20073 7650
rect 19973 7600 20073 7616
rect 5511 6323 6711 6339
rect 5511 6289 5527 6323
rect 6695 6289 6711 6323
rect 5511 6251 6711 6289
rect 5511 6013 6711 6051
rect 5511 5979 5527 6013
rect 6695 5979 6711 6013
rect 5511 5963 6711 5979
rect 7167 6323 8367 6339
rect 7167 6289 7183 6323
rect 8351 6289 8367 6323
rect 7167 6251 8367 6289
rect 7167 6013 8367 6051
rect 7167 5979 7183 6013
rect 8351 5979 8367 6013
rect 7167 5963 8367 5979
rect 16593 7115 16681 7131
rect 16593 5147 16609 7115
rect 16643 5147 16681 7115
rect 16593 5131 16681 5147
rect 16881 7115 16969 7131
rect 16881 5147 16919 7115
rect 16953 5147 16969 7115
rect 16881 5131 16969 5147
rect 17179 7115 17267 7131
rect 17179 5147 17195 7115
rect 17229 5147 17267 7115
rect 17179 5131 17267 5147
rect 17467 7115 17555 7131
rect 17467 5147 17505 7115
rect 17539 5147 17555 7115
rect 17467 5131 17555 5147
rect 17765 7115 17853 7131
rect 17765 5147 17781 7115
rect 17815 5147 17853 7115
rect 17765 5131 17853 5147
rect 18053 7115 18141 7131
rect 18053 5147 18091 7115
rect 18125 5147 18141 7115
rect 18053 5131 18141 5147
rect 16593 4653 16681 4669
rect 16593 2685 16609 4653
rect 16643 2685 16681 4653
rect 16593 2669 16681 2685
rect 16881 4653 16969 4669
rect 16881 2685 16919 4653
rect 16953 2685 16969 4653
rect 16881 2669 16969 2685
rect 17179 4653 17267 4669
rect 17179 2685 17195 4653
rect 17229 2685 17267 4653
rect 17179 2669 17267 2685
rect 17467 4653 17555 4669
rect 17467 2685 17505 4653
rect 17539 2685 17555 4653
rect 17467 2669 17555 2685
rect 17765 4653 17853 4669
rect 17765 2685 17781 4653
rect 17815 2685 17853 4653
rect 17765 2669 17853 2685
rect 18053 4653 18141 4669
rect 18053 2685 18091 4653
rect 18125 2685 18141 4653
rect 18053 2669 18141 2685
rect 21649 7883 21737 7899
rect 21649 6115 21665 7883
rect 21699 6115 21737 7883
rect 21649 6099 21737 6115
rect 23737 7883 23825 7899
rect 23737 6115 23775 7883
rect 23809 6115 23825 7883
rect 23737 6099 23825 6115
rect 24734 7883 24831 7899
rect 24734 7715 24750 7883
rect 24784 7715 24831 7883
rect 24734 7699 24831 7715
rect 25631 7883 25728 7899
rect 25631 7715 25678 7883
rect 25712 7715 25728 7883
rect 25631 7699 25728 7715
rect 21649 5633 21737 5649
rect 21649 3865 21665 5633
rect 21699 3865 21737 5633
rect 21649 3849 21737 3865
rect 23737 5633 23825 5649
rect 23737 3865 23775 5633
rect 23809 3865 23825 5633
rect 23737 3849 23825 3865
rect 24734 7177 24831 7193
rect 24734 7009 24750 7177
rect 24784 7009 24831 7177
rect 24734 6993 24831 7009
rect 26531 7177 26628 7193
rect 26531 7009 26578 7177
rect 26612 7009 26628 7177
rect 26531 6993 26628 7009
rect 24734 6919 24831 6935
rect 24734 6751 24750 6919
rect 24784 6751 24831 6919
rect 24734 6735 24831 6751
rect 26531 6919 26628 6935
rect 26531 6751 26578 6919
rect 26612 6751 26628 6919
rect 26531 6735 26628 6751
rect 24734 6661 24831 6677
rect 24734 6493 24750 6661
rect 24784 6493 24831 6661
rect 24734 6477 24831 6493
rect 26531 6661 26628 6677
rect 26531 6493 26578 6661
rect 26612 6493 26628 6661
rect 26531 6477 26628 6493
rect 24734 6403 24831 6419
rect 24734 6235 24750 6403
rect 24784 6235 24831 6403
rect 24734 6219 24831 6235
rect 26531 6403 26628 6419
rect 26531 6235 26578 6403
rect 26612 6235 26628 6403
rect 26531 6219 26628 6235
rect 24734 6145 24831 6161
rect 24734 5977 24750 6145
rect 24784 5977 24831 6145
rect 24734 5961 24831 5977
rect 26531 6145 26628 6161
rect 26531 5977 26578 6145
rect 26612 5977 26628 6145
rect 26531 5961 26628 5977
rect 24734 5887 24831 5903
rect 24734 5719 24750 5887
rect 24784 5719 24831 5887
rect 24734 5703 24831 5719
rect 26531 5887 26628 5903
rect 26531 5719 26578 5887
rect 26612 5719 26628 5887
rect 26531 5703 26628 5719
rect 24734 5629 24831 5645
rect 24734 5461 24750 5629
rect 24784 5461 24831 5629
rect 24734 5445 24831 5461
rect 26531 5629 26628 5645
rect 26531 5461 26578 5629
rect 26612 5461 26628 5629
rect 26531 5445 26628 5461
rect 24734 5371 24831 5387
rect 24734 5203 24750 5371
rect 24784 5203 24831 5371
rect 24734 5187 24831 5203
rect 26531 5371 26628 5387
rect 26531 5203 26578 5371
rect 26612 5203 26628 5371
rect 26531 5187 26628 5203
rect 21492 2999 21692 3015
rect 21492 2965 21508 2999
rect 21676 2965 21692 2999
rect 21492 2927 21692 2965
rect 21750 2999 21950 3015
rect 21750 2965 21766 2999
rect 21934 2965 21950 2999
rect 21750 2927 21950 2965
rect 22008 2999 22208 3015
rect 22008 2965 22024 2999
rect 22192 2965 22208 2999
rect 22008 2927 22208 2965
rect 22266 2999 22466 3015
rect 22266 2965 22282 2999
rect 22450 2965 22466 2999
rect 22266 2927 22466 2965
rect 22524 2999 22724 3015
rect 22524 2965 22540 2999
rect 22708 2965 22724 2999
rect 22524 2927 22724 2965
rect 22782 2999 22982 3015
rect 22782 2965 22798 2999
rect 22966 2965 22982 2999
rect 22782 2927 22982 2965
rect 23040 2999 23240 3015
rect 23040 2965 23056 2999
rect 23224 2965 23240 2999
rect 23040 2927 23240 2965
rect 23298 2999 23498 3015
rect 23298 2965 23314 2999
rect 23482 2965 23498 2999
rect 23298 2927 23498 2965
rect 23556 2999 23756 3015
rect 23556 2965 23572 2999
rect 23740 2965 23756 2999
rect 23556 2927 23756 2965
rect 23814 2999 24014 3015
rect 23814 2965 23830 2999
rect 23998 2965 24014 2999
rect 23814 2927 24014 2965
rect 21492 1889 21692 1927
rect 21492 1855 21508 1889
rect 21676 1855 21692 1889
rect 21492 1839 21692 1855
rect 21750 1889 21950 1927
rect 21750 1855 21766 1889
rect 21934 1855 21950 1889
rect 21750 1839 21950 1855
rect 22008 1889 22208 1927
rect 22008 1855 22024 1889
rect 22192 1855 22208 1889
rect 22008 1839 22208 1855
rect 22266 1889 22466 1927
rect 22266 1855 22282 1889
rect 22450 1855 22466 1889
rect 22266 1839 22466 1855
rect 22524 1889 22724 1927
rect 22524 1855 22540 1889
rect 22708 1855 22724 1889
rect 22524 1839 22724 1855
rect 22782 1889 22982 1927
rect 22782 1855 22798 1889
rect 22966 1855 22982 1889
rect 22782 1839 22982 1855
rect 23040 1889 23240 1927
rect 23040 1855 23056 1889
rect 23224 1855 23240 1889
rect 23040 1839 23240 1855
rect 23298 1889 23498 1927
rect 23298 1855 23314 1889
rect 23482 1855 23498 1889
rect 23298 1839 23498 1855
rect 23556 1889 23756 1927
rect 23556 1855 23572 1889
rect 23740 1855 23756 1889
rect 23556 1839 23756 1855
rect 23814 1889 24014 1927
rect 23814 1855 23830 1889
rect 23998 1855 24014 1889
rect 23814 1839 24014 1855
rect 24578 3775 24666 3791
rect 24578 2007 24594 3775
rect 24628 2007 24666 3775
rect 24578 1991 24666 2007
rect 26666 3775 26754 3791
rect 26666 2007 26704 3775
rect 26738 2007 26754 3775
rect 26666 1991 26754 2007
<< polycont >>
rect 6295 30965 8263 30999
rect 6295 30637 8263 30671
rect 8621 30965 10589 30999
rect 8621 30637 10589 30671
rect 6080 20072 6114 24040
rect 6290 20072 6324 24040
rect 6566 20072 6600 24040
rect 6776 20072 6810 24040
rect 7052 20072 7086 24040
rect 7262 20072 7296 24040
rect 7538 20072 7572 24040
rect 7748 20072 7782 24040
rect 8024 20072 8058 24040
rect 8234 20072 8268 24040
rect 8510 20072 8544 24040
rect 8720 20072 8754 24040
rect 8996 20072 9030 24040
rect 9206 20072 9240 24040
rect 9482 20072 9516 24040
rect 9692 20072 9726 24040
rect 9968 20072 10002 24040
rect 10178 20072 10212 24040
rect 10454 20072 10488 24040
rect 10664 20072 10698 24040
rect 11403 23257 15371 23291
rect 11403 22547 15371 22581
rect 15859 23657 19827 23691
rect 15859 22547 19827 22581
rect 11410 21985 15378 22019
rect 11410 20875 15378 20909
rect 15859 21985 19827 22019
rect 15859 21275 19827 21309
rect 6420 19098 10388 19132
rect 6420 18670 10388 18704
rect 6420 18562 10388 18596
rect 6420 18134 10388 18168
rect 6420 17698 10388 17732
rect 6420 16970 10388 17004
rect 11508 19098 15476 19132
rect 11508 16970 15476 17004
rect 15834 19098 19802 19132
rect 15834 16970 19802 17004
rect 8430 14894 10388 14928
rect 8430 14566 10388 14600
rect 11508 16694 15476 16728
rect 11508 14566 15476 14600
rect 15834 16694 19802 16728
rect 15834 14566 19802 14600
rect 20818 14738 20852 18706
rect 21046 14738 21080 18706
rect 21322 14738 21356 18706
rect 21550 14738 21584 18706
rect 8135 12370 10113 12404
rect 8135 12042 10113 12076
rect 6135 11607 10103 11641
rect 6135 11079 10103 11113
rect 6247 10621 6695 10655
rect 6247 9993 6695 10027
rect 7183 10621 7631 10655
rect 7183 9993 7631 10027
rect 9113 10639 9561 10673
rect 9113 10011 9561 10045
rect 10045 10639 10493 10673
rect 10045 10011 10493 10045
rect 12095 10912 12163 10946
rect 12253 10912 12321 10946
rect 12411 10912 12479 10946
rect 12569 10912 12637 10946
rect 12095 10584 12163 10618
rect 12253 10584 12321 10618
rect 12411 10584 12479 10618
rect 12569 10584 12637 10618
rect 6247 9579 6695 9613
rect 6247 8951 6695 8985
rect 7183 9579 7631 9613
rect 7183 8951 7631 8985
rect 9113 9554 9561 9588
rect 9113 8926 9561 8960
rect 10045 9554 10493 9588
rect 10045 8926 10493 8960
rect 11479 9688 11547 9722
rect 11479 9378 11547 9412
rect 12035 9688 12103 9722
rect 12035 9378 12103 9412
rect 12591 9688 12659 9722
rect 12591 9378 12659 9412
rect 13147 9688 13215 9722
rect 13147 9378 13215 9412
rect 5527 8437 6695 8471
rect 5527 8127 6695 8161
rect 7183 8437 8351 8471
rect 7183 8127 8351 8161
rect 9113 8437 9521 8471
rect 9113 8127 9521 8161
rect 10085 8438 10493 8472
rect 10085 8128 10493 8162
rect 5527 7721 6695 7755
rect 5527 7411 6695 7445
rect 7183 7721 8351 7755
rect 7183 7411 8351 7445
rect 5527 7005 6695 7039
rect 5527 6695 6695 6729
rect 7183 7005 8351 7039
rect 7183 6695 8351 6729
rect 16671 9726 16739 9760
rect 16829 9726 16897 9760
rect 16987 9726 17055 9760
rect 17145 9726 17213 9760
rect 17303 9726 17371 9760
rect 17461 9726 17529 9760
rect 17619 9726 17687 9760
rect 17777 9726 17845 9760
rect 17935 9726 18003 9760
rect 18093 9726 18161 9760
rect 18251 9726 18319 9760
rect 18409 9726 18477 9760
rect 18567 9726 18635 9760
rect 18725 9726 18793 9760
rect 18883 9726 18951 9760
rect 19041 9726 19109 9760
rect 19199 9726 19267 9760
rect 19357 9726 19425 9760
rect 19515 9726 19583 9760
rect 19673 9726 19741 9760
rect 19831 9726 19899 9760
rect 19989 9726 20057 9760
rect 16671 7616 16739 7650
rect 16829 7616 16897 7650
rect 16987 7616 17055 7650
rect 17145 7616 17213 7650
rect 17303 7616 17371 7650
rect 17461 7616 17529 7650
rect 17619 7616 17687 7650
rect 17777 7616 17845 7650
rect 17935 7616 18003 7650
rect 18093 7616 18161 7650
rect 18251 7616 18319 7650
rect 18409 7616 18477 7650
rect 18567 7616 18635 7650
rect 18725 7616 18793 7650
rect 18883 7616 18951 7650
rect 19041 7616 19109 7650
rect 19199 7616 19267 7650
rect 19357 7616 19425 7650
rect 19515 7616 19583 7650
rect 19673 7616 19741 7650
rect 19831 7616 19899 7650
rect 19989 7616 20057 7650
rect 5527 6289 6695 6323
rect 5527 5979 6695 6013
rect 7183 6289 8351 6323
rect 7183 5979 8351 6013
rect 16609 5147 16643 7115
rect 16919 5147 16953 7115
rect 17195 5147 17229 7115
rect 17505 5147 17539 7115
rect 17781 5147 17815 7115
rect 18091 5147 18125 7115
rect 16609 2685 16643 4653
rect 16919 2685 16953 4653
rect 17195 2685 17229 4653
rect 17505 2685 17539 4653
rect 17781 2685 17815 4653
rect 18091 2685 18125 4653
rect 21665 6115 21699 7883
rect 23775 6115 23809 7883
rect 24750 7715 24784 7883
rect 25678 7715 25712 7883
rect 21665 3865 21699 5633
rect 23775 3865 23809 5633
rect 24750 7009 24784 7177
rect 26578 7009 26612 7177
rect 24750 6751 24784 6919
rect 26578 6751 26612 6919
rect 24750 6493 24784 6661
rect 26578 6493 26612 6661
rect 24750 6235 24784 6403
rect 26578 6235 26612 6403
rect 24750 5977 24784 6145
rect 26578 5977 26612 6145
rect 24750 5719 24784 5887
rect 26578 5719 26612 5887
rect 24750 5461 24784 5629
rect 26578 5461 26612 5629
rect 24750 5203 24784 5371
rect 26578 5203 26612 5371
rect 21508 2965 21676 2999
rect 21766 2965 21934 2999
rect 22024 2965 22192 2999
rect 22282 2965 22450 2999
rect 22540 2965 22708 2999
rect 22798 2965 22966 2999
rect 23056 2965 23224 2999
rect 23314 2965 23482 2999
rect 23572 2965 23740 2999
rect 23830 2965 23998 2999
rect 21508 1855 21676 1889
rect 21766 1855 21934 1889
rect 22024 1855 22192 1889
rect 22282 1855 22450 1889
rect 22540 1855 22708 1889
rect 22798 1855 22966 1889
rect 23056 1855 23224 1889
rect 23314 1855 23482 1889
rect 23572 1855 23740 1889
rect 23830 1855 23998 1889
rect 24594 2007 24628 3775
rect 26704 2007 26738 3775
<< xpolycontact >>
rect 2786 41806 2856 42238
rect 2786 36406 2856 36838
rect 3082 41806 3152 42238
rect 3082 36406 3152 36838
rect 3378 41806 3448 42238
rect 3378 36406 3448 36838
rect 3674 41806 3744 42238
rect 3674 36406 3744 36838
rect 3970 41806 4040 42238
rect 3970 36406 4040 36838
rect 4266 41806 4336 42238
rect 4266 36406 4336 36838
rect 4562 41806 4632 42238
rect 4562 36406 4632 36838
rect 4858 41806 4928 42238
rect 4858 36406 4928 36838
rect 5154 41806 5224 42238
rect 5154 36406 5224 36838
rect 5450 41806 5520 42238
rect 5450 36406 5520 36838
rect 2786 35748 2856 36180
rect 2786 30348 2856 30780
rect 3082 35748 3152 36180
rect 3082 30348 3152 30780
rect 3378 35748 3448 36180
rect 3378 30348 3448 30780
rect 3674 35748 3744 36180
rect 3674 30348 3744 30780
rect 3970 35748 4040 36180
rect 3970 30348 4040 30780
rect 4266 35748 4336 36180
rect 4266 30348 4336 30780
rect 4562 35748 4632 36180
rect 4562 30348 4632 30780
rect 4858 35748 4928 36180
rect 4858 30348 4928 30780
rect 5154 35748 5224 36180
rect 5154 30348 5224 30780
rect 5450 35748 5520 36180
rect 5450 30348 5520 30780
rect 7586 28043 8018 28113
rect 9886 28043 10318 28113
rect 10544 28043 10976 28113
rect 12844 28043 13276 28113
rect 7586 27747 8018 27817
rect 9886 27747 10318 27817
rect 10544 27747 10976 27817
rect 12844 27747 13276 27817
rect 7586 27451 8018 27521
rect 9886 27451 10318 27521
rect 10544 27451 10976 27521
rect 12844 27451 13276 27521
rect 7586 27155 8018 27225
rect 9886 27155 10318 27225
rect 10544 27155 10976 27225
rect 12844 27155 13276 27225
rect 7586 26859 8018 26929
rect 9886 26859 10318 26929
rect 10544 26859 10976 26929
rect 12844 26859 13276 26929
rect 7586 26563 8018 26633
rect 9886 26563 10318 26633
rect 10544 26563 10976 26633
rect 12844 26563 13276 26633
rect 7586 26267 8018 26337
rect 9886 26267 10318 26337
rect 10544 26267 10976 26337
rect 12844 26267 13276 26337
rect 7586 25971 8018 26041
rect 9886 25971 10318 26041
rect 10544 25971 10976 26041
rect 12844 25971 13276 26041
rect 7586 25675 8018 25745
rect 9886 25675 10318 25745
rect 10544 25675 10976 25745
rect 12844 25675 13276 25745
rect 7586 25379 8018 25449
rect 9886 25379 10318 25449
rect 10544 25379 10976 25449
rect 12844 25379 13276 25449
rect 7586 25083 8018 25153
rect 9886 25083 10318 25153
rect 10544 25083 10976 25153
rect 12844 25083 13276 25153
rect 7586 24787 8018 24857
rect 9886 24787 10318 24857
rect 10544 24787 10976 24857
rect 12844 24787 13276 24857
rect 14097 10265 14167 10697
rect 14097 6765 14167 7197
rect 14393 10265 14463 10697
rect 14393 6765 14463 7197
rect 14689 10265 14759 10697
rect 14689 6765 14759 7197
rect 14985 10265 15055 10697
rect 14985 6765 15055 7197
rect 15281 10265 15351 10697
rect 15281 6765 15351 7197
rect 15577 10265 15647 10697
rect 15577 6765 15647 7197
rect 15873 10265 15943 10697
rect 15873 6765 15943 7197
rect 16169 10265 16239 10697
rect 16169 6765 16239 7197
rect 14097 6107 14167 6539
rect 14097 2607 14167 3039
rect 14393 6107 14463 6539
rect 14393 2607 14463 3039
rect 14689 6107 14759 6539
rect 14689 2607 14759 3039
rect 14985 6107 15055 6539
rect 14985 2607 15055 3039
rect 15281 6107 15351 6539
rect 15281 2607 15351 3039
rect 15577 6107 15647 6539
rect 15577 2607 15647 3039
rect 15873 6107 15943 6539
rect 15873 2607 15943 3039
rect 16169 6107 16239 6539
rect 16169 2607 16239 3039
rect 18714 5807 18784 6239
rect 18714 2607 18784 3039
rect 19010 5807 19080 6239
rect 19010 2607 19080 3039
rect 19306 5807 19376 6239
rect 19306 2607 19376 3039
rect 19602 5807 19672 6239
rect 19602 2607 19672 3039
<< xpolyres >>
rect 2786 36838 2856 41806
rect 3082 36838 3152 41806
rect 3378 36838 3448 41806
rect 3674 36838 3744 41806
rect 3970 36838 4040 41806
rect 4266 36838 4336 41806
rect 4562 36838 4632 41806
rect 4858 36838 4928 41806
rect 5154 36838 5224 41806
rect 5450 36838 5520 41806
rect 2786 30780 2856 35748
rect 3082 30780 3152 35748
rect 3378 30780 3448 35748
rect 3674 30780 3744 35748
rect 3970 30780 4040 35748
rect 4266 30780 4336 35748
rect 4562 30780 4632 35748
rect 4858 30780 4928 35748
rect 5154 30780 5224 35748
rect 5450 30780 5520 35748
rect 8018 28043 9886 28113
rect 10976 28043 12844 28113
rect 8018 27747 9886 27817
rect 10976 27747 12844 27817
rect 8018 27451 9886 27521
rect 10976 27451 12844 27521
rect 8018 27155 9886 27225
rect 10976 27155 12844 27225
rect 8018 26859 9886 26929
rect 10976 26859 12844 26929
rect 8018 26563 9886 26633
rect 10976 26563 12844 26633
rect 8018 26267 9886 26337
rect 10976 26267 12844 26337
rect 8018 25971 9886 26041
rect 10976 25971 12844 26041
rect 8018 25675 9886 25745
rect 10976 25675 12844 25745
rect 8018 25379 9886 25449
rect 10976 25379 12844 25449
rect 8018 25083 9886 25153
rect 10976 25083 12844 25153
rect 8018 24787 9886 24857
rect 10976 24787 12844 24857
rect 14097 7197 14167 10265
rect 14393 7197 14463 10265
rect 14689 7197 14759 10265
rect 14985 7197 15055 10265
rect 15281 7197 15351 10265
rect 15577 7197 15647 10265
rect 15873 7197 15943 10265
rect 16169 7197 16239 10265
rect 14097 3039 14167 6107
rect 14393 3039 14463 6107
rect 14689 3039 14759 6107
rect 14985 3039 15055 6107
rect 15281 3039 15351 6107
rect 15577 3039 15647 6107
rect 15873 3039 15943 6107
rect 16169 3039 16239 6107
rect 18714 3039 18784 5807
rect 19010 3039 19080 5807
rect 19306 3039 19376 5807
rect 19602 3039 19672 5807
<< locali >>
rect 2405 42620 5794 42622
rect 2405 42578 5841 42620
rect 2405 42577 2669 42578
rect 2405 30063 2431 42577
rect 5829 42347 5841 42578
rect 2681 42334 2752 42347
rect 2890 42334 3048 42347
rect 3186 42334 3344 42347
rect 3482 42334 3640 42347
rect 3778 42334 3936 42347
rect 4074 42334 4232 42347
rect 4370 42334 4528 42347
rect 4666 42334 4824 42347
rect 4962 42334 5120 42347
rect 5258 42334 5416 42347
rect 5554 42334 5613 42347
rect 2681 42311 5613 42334
rect 2681 42272 2716 42311
rect 2690 36372 2716 42272
rect 2952 42272 2986 42311
rect 2681 36310 2716 36372
rect 3248 42272 3282 42311
rect 2952 36310 2986 36372
rect 3544 42272 3578 42311
rect 3248 36310 3282 36372
rect 3840 42272 3874 42311
rect 3544 36310 3578 36372
rect 4136 42272 4170 42311
rect 3840 36310 3874 36372
rect 4432 42272 4466 42311
rect 4136 36310 4170 36372
rect 4728 42272 4762 42311
rect 4432 36310 4466 36372
rect 5024 42272 5058 42311
rect 4728 36310 4762 36372
rect 5320 42272 5354 42311
rect 5024 36310 5058 36372
rect 5320 36310 5354 36372
rect 5590 36310 5613 42311
rect 2681 36276 2752 36310
rect 2890 36276 3048 36310
rect 3186 36276 3344 36310
rect 3482 36276 3640 36310
rect 3778 36276 3936 36310
rect 4074 36276 4232 36310
rect 4370 36276 4528 36310
rect 4666 36276 4824 36310
rect 4962 36276 5120 36310
rect 5258 36276 5416 36310
rect 5554 36276 5613 36310
rect 2681 36214 2716 36276
rect 2690 30314 2716 36214
rect 2952 36214 2986 36276
rect 2681 30294 2716 30314
rect 3248 36214 3282 36276
rect 2952 30294 2986 30314
rect 3544 36214 3578 36276
rect 3248 30294 3282 30314
rect 3840 36214 3874 36276
rect 3544 30294 3578 30314
rect 4136 36214 4170 36276
rect 3840 30294 3874 30314
rect 4432 36214 4466 36276
rect 4136 30294 4170 30314
rect 4728 36214 4762 36276
rect 4432 30294 4466 30314
rect 5024 36214 5058 36276
rect 4728 30294 4762 30314
rect 5320 36214 5354 36276
rect 5024 30294 5058 30314
rect 5320 30294 5354 30314
rect 5590 30294 5613 36276
rect 2681 30252 5613 30294
rect 2681 30245 2752 30252
rect 2890 30245 3048 30252
rect 3186 30245 3344 30252
rect 3482 30245 3640 30252
rect 3778 30245 3936 30252
rect 4074 30245 4232 30252
rect 4370 30245 4528 30252
rect 4666 30245 4824 30252
rect 4962 30245 5120 30252
rect 5258 30245 5416 30252
rect 5554 30245 5613 30252
rect 2405 30058 2491 30063
rect 5815 30058 5841 42347
rect 6022 31147 6032 31284
rect 6022 30450 6028 31147
rect 10883 31118 10904 31284
rect 6143 31103 6195 31118
rect 8363 31103 8521 31118
rect 10689 31103 10759 31118
rect 6143 31098 10759 31103
rect 6143 30547 6160 31098
rect 8425 31041 8459 31098
rect 6279 30965 6295 30999
rect 8263 30965 8279 30999
rect 6233 30906 6267 30922
rect 6233 30714 6267 30730
rect 8291 30906 8325 30922
rect 8291 30714 8325 30730
rect 6279 30637 6295 30671
rect 8263 30637 8279 30671
rect 10748 31041 10759 31098
rect 8605 30965 8621 30999
rect 10589 30965 10605 30999
rect 8559 30906 8593 30922
rect 8559 30714 8593 30730
rect 10617 30906 10651 30922
rect 10617 30714 10651 30730
rect 8605 30637 8621 30671
rect 10589 30637 10605 30671
rect 8425 30547 8459 30595
rect 10748 30595 10751 31041
rect 10748 30547 10759 30595
rect 6143 30536 10759 30547
rect 10874 30536 10904 31118
rect 6022 30351 6031 30450
rect 10882 30351 10904 30536
rect 6022 30335 10904 30351
rect 2405 30028 5841 30058
rect 7335 28343 17633 28357
rect 7335 28190 7370 28343
rect 17591 28190 17633 28343
rect 7335 24690 7371 28190
rect 7490 28183 13405 28190
rect 7490 27974 7495 28183
rect 10377 28147 10475 28183
rect 10377 28009 10414 28147
rect 10448 28009 10475 28147
rect 13370 28147 13405 28183
rect 17590 28183 17633 28190
rect 10377 27974 10475 28009
rect 13370 28009 13372 28147
rect 13844 28046 13921 28050
rect 13955 28046 14011 28050
rect 14045 28046 14101 28050
rect 14135 28046 14191 28050
rect 14225 28046 14281 28050
rect 14315 28046 14371 28050
rect 14405 28046 14461 28050
rect 14495 28046 14551 28050
rect 14585 28046 14641 28050
rect 14675 28046 14739 28050
rect 13844 28027 14739 28046
rect 13370 27974 13405 28009
rect 13844 27986 13882 28027
rect 7490 27947 13405 27974
rect 7490 27913 7552 27947
rect 10352 27913 10510 27947
rect 13310 27913 13405 27947
rect 13863 27952 13882 27986
rect 14700 27967 14739 28027
rect 15181 28046 15265 28050
rect 15299 28046 15355 28050
rect 15389 28046 15445 28050
rect 15479 28046 15535 28050
rect 15569 28046 15625 28050
rect 15659 28046 15715 28050
rect 15749 28046 15805 28050
rect 15839 28046 15895 28050
rect 15929 28046 15985 28050
rect 16019 28046 16084 28050
rect 15181 28027 16084 28046
rect 15181 27986 15226 28027
rect 7490 27863 13405 27913
rect 13844 27896 13882 27952
rect 7490 27681 7495 27863
rect 10377 27851 10475 27863
rect 10377 27713 10414 27851
rect 10448 27713 10475 27851
rect 13370 27851 13405 27863
rect 10377 27681 10475 27713
rect 13370 27713 13372 27851
rect 13863 27862 13882 27896
rect 13844 27806 13882 27862
rect 13863 27772 13882 27806
rect 13844 27716 13882 27772
rect 13370 27681 13405 27713
rect 7490 27651 13405 27681
rect 13863 27682 13882 27716
rect 7490 27617 7552 27651
rect 10352 27617 10510 27651
rect 13310 27617 13405 27651
rect 13844 27626 13882 27682
rect 7490 27570 13405 27617
rect 13863 27592 13882 27626
rect 7490 27387 7495 27570
rect 10377 27555 10475 27570
rect 10377 27417 10414 27555
rect 10448 27417 10475 27555
rect 13370 27555 13405 27570
rect 10377 27387 10475 27417
rect 13370 27417 13372 27555
rect 13844 27536 13882 27592
rect 13863 27502 13882 27536
rect 13844 27446 13882 27502
rect 13370 27387 13405 27417
rect 13863 27412 13882 27446
rect 7490 27355 13405 27387
rect 13844 27356 13882 27412
rect 7490 27321 7552 27355
rect 10352 27321 10510 27355
rect 13310 27321 13405 27355
rect 7490 27276 13405 27321
rect 13863 27322 13882 27356
rect 7490 27094 7495 27276
rect 10377 27259 10475 27276
rect 10377 27121 10414 27259
rect 10448 27121 10475 27259
rect 13370 27259 13405 27276
rect 13844 27266 13882 27322
rect 13944 27904 14638 27965
rect 13944 27870 14003 27904
rect 14037 27892 14093 27904
rect 14065 27870 14093 27892
rect 14127 27892 14183 27904
rect 14127 27870 14131 27892
rect 13944 27858 14031 27870
rect 14065 27858 14131 27870
rect 14165 27870 14183 27892
rect 14217 27892 14273 27904
rect 14217 27870 14231 27892
rect 14165 27858 14231 27870
rect 14265 27870 14273 27892
rect 14307 27892 14363 27904
rect 14397 27892 14453 27904
rect 14487 27892 14543 27904
rect 14307 27870 14331 27892
rect 14397 27870 14431 27892
rect 14487 27870 14531 27892
rect 14577 27870 14638 27904
rect 14265 27858 14331 27870
rect 14365 27858 14431 27870
rect 14465 27858 14531 27870
rect 14565 27858 14638 27870
rect 13944 27814 14638 27858
rect 13944 27780 14003 27814
rect 14037 27792 14093 27814
rect 14065 27780 14093 27792
rect 14127 27792 14183 27814
rect 14127 27780 14131 27792
rect 13944 27758 14031 27780
rect 14065 27758 14131 27780
rect 14165 27780 14183 27792
rect 14217 27792 14273 27814
rect 14217 27780 14231 27792
rect 14165 27758 14231 27780
rect 14265 27780 14273 27792
rect 14307 27792 14363 27814
rect 14397 27792 14453 27814
rect 14487 27792 14543 27814
rect 14307 27780 14331 27792
rect 14397 27780 14431 27792
rect 14487 27780 14531 27792
rect 14577 27780 14638 27814
rect 14265 27758 14331 27780
rect 14365 27758 14431 27780
rect 14465 27758 14531 27780
rect 14565 27758 14638 27780
rect 13944 27724 14638 27758
rect 13944 27690 14003 27724
rect 14037 27692 14093 27724
rect 14065 27690 14093 27692
rect 14127 27692 14183 27724
rect 14127 27690 14131 27692
rect 13944 27658 14031 27690
rect 14065 27658 14131 27690
rect 14165 27690 14183 27692
rect 14217 27692 14273 27724
rect 14217 27690 14231 27692
rect 14165 27658 14231 27690
rect 14265 27690 14273 27692
rect 14307 27692 14363 27724
rect 14397 27692 14453 27724
rect 14487 27692 14543 27724
rect 14307 27690 14331 27692
rect 14397 27690 14431 27692
rect 14487 27690 14531 27692
rect 14577 27690 14638 27724
rect 14265 27658 14331 27690
rect 14365 27658 14431 27690
rect 14465 27658 14531 27690
rect 14565 27658 14638 27690
rect 13944 27634 14638 27658
rect 13944 27600 14003 27634
rect 14037 27600 14093 27634
rect 14127 27600 14183 27634
rect 14217 27600 14273 27634
rect 14307 27600 14363 27634
rect 14397 27600 14453 27634
rect 14487 27600 14543 27634
rect 14577 27600 14638 27634
rect 13944 27592 14638 27600
rect 13944 27558 14031 27592
rect 14065 27558 14131 27592
rect 14165 27558 14231 27592
rect 14265 27558 14331 27592
rect 14365 27558 14431 27592
rect 14465 27558 14531 27592
rect 14565 27558 14638 27592
rect 13944 27544 14638 27558
rect 13944 27510 14003 27544
rect 14037 27510 14093 27544
rect 14127 27510 14183 27544
rect 14217 27510 14273 27544
rect 14307 27510 14363 27544
rect 14397 27510 14453 27544
rect 14487 27510 14543 27544
rect 14577 27510 14638 27544
rect 13944 27492 14638 27510
rect 13944 27458 14031 27492
rect 14065 27458 14131 27492
rect 14165 27458 14231 27492
rect 14265 27458 14331 27492
rect 14365 27458 14431 27492
rect 14465 27458 14531 27492
rect 14565 27458 14638 27492
rect 13944 27454 14638 27458
rect 13944 27420 14003 27454
rect 14037 27420 14093 27454
rect 14127 27420 14183 27454
rect 14217 27420 14273 27454
rect 14307 27420 14363 27454
rect 14397 27420 14453 27454
rect 14487 27420 14543 27454
rect 14577 27420 14638 27454
rect 13944 27392 14638 27420
rect 13944 27364 14031 27392
rect 14065 27364 14131 27392
rect 13944 27330 14003 27364
rect 14065 27358 14093 27364
rect 14037 27330 14093 27358
rect 14127 27358 14131 27364
rect 14165 27364 14231 27392
rect 14165 27358 14183 27364
rect 14127 27330 14183 27358
rect 14217 27358 14231 27364
rect 14265 27364 14331 27392
rect 14365 27364 14431 27392
rect 14465 27364 14531 27392
rect 14565 27364 14638 27392
rect 14265 27358 14273 27364
rect 14217 27330 14273 27358
rect 14307 27358 14331 27364
rect 14397 27358 14431 27364
rect 14487 27358 14531 27364
rect 14307 27330 14363 27358
rect 14397 27330 14453 27358
rect 14487 27330 14543 27358
rect 14577 27330 14638 27364
rect 13944 27271 14638 27330
rect 14700 27933 14719 27967
rect 14700 27877 14739 27933
rect 15207 27952 15226 27986
rect 16044 27967 16084 28027
rect 16526 28046 16609 28050
rect 16643 28046 16699 28050
rect 16733 28046 16789 28050
rect 16823 28046 16879 28050
rect 16913 28046 16969 28050
rect 17003 28046 17059 28050
rect 17093 28046 17149 28050
rect 17183 28046 17239 28050
rect 17273 28046 17329 28050
rect 17363 28046 17424 28050
rect 16526 28027 17424 28046
rect 16526 27986 16570 28027
rect 15181 27896 15226 27952
rect 14700 27843 14719 27877
rect 14700 27825 14739 27843
rect 15207 27862 15226 27896
rect 15181 27825 15226 27862
rect 14700 27806 15226 27825
rect 14700 27787 15173 27806
rect 14700 27753 14719 27787
rect 14753 27786 15173 27787
rect 14753 27753 14867 27786
rect 14700 27752 14867 27753
rect 14901 27752 15024 27786
rect 15058 27772 15173 27786
rect 15207 27772 15226 27806
rect 15058 27752 15226 27772
rect 14700 27716 15226 27752
rect 14700 27697 15173 27716
rect 14700 27663 14719 27697
rect 14753 27696 15173 27697
rect 14753 27663 14867 27696
rect 14700 27662 14867 27663
rect 14901 27662 15024 27696
rect 15058 27682 15173 27696
rect 15207 27682 15226 27716
rect 15058 27662 15226 27682
rect 14700 27626 15226 27662
rect 14700 27607 15173 27626
rect 14700 27573 14719 27607
rect 14753 27606 15173 27607
rect 14753 27573 14867 27606
rect 14700 27572 14867 27573
rect 14901 27572 15024 27606
rect 15058 27592 15173 27606
rect 15207 27592 15226 27626
rect 15058 27572 15226 27592
rect 14700 27536 15226 27572
rect 14700 27517 15173 27536
rect 14700 27483 14719 27517
rect 14753 27516 15173 27517
rect 14753 27483 14867 27516
rect 14700 27482 14867 27483
rect 14901 27482 15024 27516
rect 15058 27502 15173 27516
rect 15207 27502 15226 27536
rect 15058 27482 15226 27502
rect 14700 27446 15226 27482
rect 14700 27427 15173 27446
rect 14700 27393 14719 27427
rect 14753 27426 15173 27427
rect 14753 27393 14867 27426
rect 14700 27392 14867 27393
rect 14901 27392 15024 27426
rect 15058 27412 15173 27426
rect 15207 27412 15226 27446
rect 15058 27392 15226 27412
rect 14700 27372 15226 27392
rect 14700 27337 14762 27372
rect 15178 27356 15226 27372
rect 14700 27303 14719 27337
rect 14753 27303 14762 27337
rect 10377 27094 10475 27121
rect 13370 27121 13372 27259
rect 13863 27232 13882 27266
rect 13844 27209 13882 27232
rect 14700 27247 14762 27303
rect 15207 27322 15226 27356
rect 15178 27266 15226 27322
rect 15288 27904 15982 27965
rect 15288 27870 15347 27904
rect 15381 27892 15437 27904
rect 15409 27870 15437 27892
rect 15471 27892 15527 27904
rect 15471 27870 15475 27892
rect 15288 27858 15375 27870
rect 15409 27858 15475 27870
rect 15509 27870 15527 27892
rect 15561 27892 15617 27904
rect 15561 27870 15575 27892
rect 15509 27858 15575 27870
rect 15609 27870 15617 27892
rect 15651 27892 15707 27904
rect 15741 27892 15797 27904
rect 15831 27892 15887 27904
rect 15651 27870 15675 27892
rect 15741 27870 15775 27892
rect 15831 27870 15875 27892
rect 15921 27870 15982 27904
rect 15609 27858 15675 27870
rect 15709 27858 15775 27870
rect 15809 27858 15875 27870
rect 15909 27858 15982 27870
rect 15288 27814 15982 27858
rect 15288 27780 15347 27814
rect 15381 27792 15437 27814
rect 15409 27780 15437 27792
rect 15471 27792 15527 27814
rect 15471 27780 15475 27792
rect 15288 27758 15375 27780
rect 15409 27758 15475 27780
rect 15509 27780 15527 27792
rect 15561 27792 15617 27814
rect 15561 27780 15575 27792
rect 15509 27758 15575 27780
rect 15609 27780 15617 27792
rect 15651 27792 15707 27814
rect 15741 27792 15797 27814
rect 15831 27792 15887 27814
rect 15651 27780 15675 27792
rect 15741 27780 15775 27792
rect 15831 27780 15875 27792
rect 15921 27780 15982 27814
rect 15609 27758 15675 27780
rect 15709 27758 15775 27780
rect 15809 27758 15875 27780
rect 15909 27758 15982 27780
rect 15288 27724 15982 27758
rect 15288 27690 15347 27724
rect 15381 27692 15437 27724
rect 15409 27690 15437 27692
rect 15471 27692 15527 27724
rect 15471 27690 15475 27692
rect 15288 27658 15375 27690
rect 15409 27658 15475 27690
rect 15509 27690 15527 27692
rect 15561 27692 15617 27724
rect 15561 27690 15575 27692
rect 15509 27658 15575 27690
rect 15609 27690 15617 27692
rect 15651 27692 15707 27724
rect 15741 27692 15797 27724
rect 15831 27692 15887 27724
rect 15651 27690 15675 27692
rect 15741 27690 15775 27692
rect 15831 27690 15875 27692
rect 15921 27690 15982 27724
rect 15609 27658 15675 27690
rect 15709 27658 15775 27690
rect 15809 27658 15875 27690
rect 15909 27658 15982 27690
rect 15288 27634 15982 27658
rect 15288 27600 15347 27634
rect 15381 27600 15437 27634
rect 15471 27600 15527 27634
rect 15561 27600 15617 27634
rect 15651 27600 15707 27634
rect 15741 27600 15797 27634
rect 15831 27600 15887 27634
rect 15921 27600 15982 27634
rect 15288 27592 15982 27600
rect 15288 27558 15375 27592
rect 15409 27558 15475 27592
rect 15509 27558 15575 27592
rect 15609 27558 15675 27592
rect 15709 27558 15775 27592
rect 15809 27558 15875 27592
rect 15909 27558 15982 27592
rect 15288 27544 15982 27558
rect 15288 27510 15347 27544
rect 15381 27510 15437 27544
rect 15471 27510 15527 27544
rect 15561 27510 15617 27544
rect 15651 27510 15707 27544
rect 15741 27510 15797 27544
rect 15831 27510 15887 27544
rect 15921 27510 15982 27544
rect 15288 27492 15982 27510
rect 15288 27458 15375 27492
rect 15409 27458 15475 27492
rect 15509 27458 15575 27492
rect 15609 27458 15675 27492
rect 15709 27458 15775 27492
rect 15809 27458 15875 27492
rect 15909 27458 15982 27492
rect 15288 27454 15982 27458
rect 15288 27420 15347 27454
rect 15381 27420 15437 27454
rect 15471 27420 15527 27454
rect 15561 27420 15617 27454
rect 15651 27420 15707 27454
rect 15741 27420 15797 27454
rect 15831 27420 15887 27454
rect 15921 27420 15982 27454
rect 15288 27392 15982 27420
rect 15288 27364 15375 27392
rect 15409 27364 15475 27392
rect 15288 27330 15347 27364
rect 15409 27358 15437 27364
rect 15381 27330 15437 27358
rect 15471 27358 15475 27364
rect 15509 27364 15575 27392
rect 15509 27358 15527 27364
rect 15471 27330 15527 27358
rect 15561 27358 15575 27364
rect 15609 27364 15675 27392
rect 15709 27364 15775 27392
rect 15809 27364 15875 27392
rect 15909 27364 15982 27392
rect 15609 27358 15617 27364
rect 15561 27330 15617 27358
rect 15651 27358 15675 27364
rect 15741 27358 15775 27364
rect 15831 27358 15875 27364
rect 15651 27330 15707 27358
rect 15741 27330 15797 27358
rect 15831 27330 15887 27358
rect 15921 27330 15982 27364
rect 15288 27271 15982 27330
rect 16044 27933 16063 27967
rect 16044 27877 16084 27933
rect 16551 27952 16570 27986
rect 17388 27967 17424 28027
rect 16526 27896 16570 27952
rect 16044 27843 16063 27877
rect 16044 27814 16084 27843
rect 16551 27862 16570 27896
rect 16526 27814 16570 27862
rect 16044 27806 16570 27814
rect 16044 27787 16517 27806
rect 16044 27753 16063 27787
rect 16097 27786 16517 27787
rect 16097 27753 16211 27786
rect 16044 27752 16211 27753
rect 16245 27752 16368 27786
rect 16402 27772 16517 27786
rect 16551 27772 16570 27806
rect 16402 27752 16570 27772
rect 16044 27716 16570 27752
rect 16044 27697 16517 27716
rect 16044 27663 16063 27697
rect 16097 27696 16517 27697
rect 16097 27663 16211 27696
rect 16044 27662 16211 27663
rect 16245 27662 16368 27696
rect 16402 27682 16517 27696
rect 16551 27682 16570 27716
rect 16402 27662 16570 27682
rect 16044 27626 16570 27662
rect 16044 27607 16517 27626
rect 16044 27573 16063 27607
rect 16097 27606 16517 27607
rect 16097 27573 16211 27606
rect 16044 27572 16211 27573
rect 16245 27572 16368 27606
rect 16402 27592 16517 27606
rect 16551 27592 16570 27626
rect 16402 27572 16570 27592
rect 16044 27536 16570 27572
rect 16044 27517 16517 27536
rect 16044 27483 16063 27517
rect 16097 27516 16517 27517
rect 16097 27483 16211 27516
rect 16044 27482 16211 27483
rect 16245 27482 16368 27516
rect 16402 27502 16517 27516
rect 16551 27502 16570 27536
rect 16402 27482 16570 27502
rect 16044 27446 16570 27482
rect 16044 27427 16517 27446
rect 16044 27393 16063 27427
rect 16097 27426 16517 27427
rect 16097 27393 16211 27426
rect 16044 27392 16211 27393
rect 16245 27392 16368 27426
rect 16402 27412 16517 27426
rect 16551 27412 16570 27446
rect 16402 27392 16570 27412
rect 16044 27372 16570 27392
rect 16044 27337 16092 27372
rect 16508 27356 16570 27372
rect 16044 27303 16063 27337
rect 14700 27213 14719 27247
rect 14753 27213 14762 27247
rect 14700 27209 14762 27213
rect 15207 27232 15226 27266
rect 13844 27190 14762 27209
rect 13844 27172 13887 27190
rect 13921 27172 13977 27190
rect 14011 27172 14067 27190
rect 14101 27156 14157 27190
rect 14191 27156 14247 27190
rect 14281 27156 14337 27190
rect 14371 27156 14427 27190
rect 14461 27156 14517 27190
rect 14551 27175 14607 27190
rect 14641 27175 14762 27190
rect 15178 27209 15226 27232
rect 16044 27247 16092 27303
rect 16508 27322 16517 27356
rect 16551 27322 16570 27356
rect 16508 27266 16570 27322
rect 16632 27904 17326 27965
rect 16632 27870 16691 27904
rect 16725 27892 16781 27904
rect 16753 27870 16781 27892
rect 16815 27892 16871 27904
rect 16815 27870 16819 27892
rect 16632 27858 16719 27870
rect 16753 27858 16819 27870
rect 16853 27870 16871 27892
rect 16905 27892 16961 27904
rect 16905 27870 16919 27892
rect 16853 27858 16919 27870
rect 16953 27870 16961 27892
rect 16995 27892 17051 27904
rect 17085 27892 17141 27904
rect 17175 27892 17231 27904
rect 16995 27870 17019 27892
rect 17085 27870 17119 27892
rect 17175 27870 17219 27892
rect 17265 27870 17326 27904
rect 16953 27858 17019 27870
rect 17053 27858 17119 27870
rect 17153 27858 17219 27870
rect 17253 27858 17326 27870
rect 16632 27814 17326 27858
rect 16632 27780 16691 27814
rect 16725 27792 16781 27814
rect 16753 27780 16781 27792
rect 16815 27792 16871 27814
rect 16815 27780 16819 27792
rect 16632 27758 16719 27780
rect 16753 27758 16819 27780
rect 16853 27780 16871 27792
rect 16905 27792 16961 27814
rect 16905 27780 16919 27792
rect 16853 27758 16919 27780
rect 16953 27780 16961 27792
rect 16995 27792 17051 27814
rect 17085 27792 17141 27814
rect 17175 27792 17231 27814
rect 16995 27780 17019 27792
rect 17085 27780 17119 27792
rect 17175 27780 17219 27792
rect 17265 27780 17326 27814
rect 16953 27758 17019 27780
rect 17053 27758 17119 27780
rect 17153 27758 17219 27780
rect 17253 27758 17326 27780
rect 16632 27724 17326 27758
rect 16632 27690 16691 27724
rect 16725 27692 16781 27724
rect 16753 27690 16781 27692
rect 16815 27692 16871 27724
rect 16815 27690 16819 27692
rect 16632 27658 16719 27690
rect 16753 27658 16819 27690
rect 16853 27690 16871 27692
rect 16905 27692 16961 27724
rect 16905 27690 16919 27692
rect 16853 27658 16919 27690
rect 16953 27690 16961 27692
rect 16995 27692 17051 27724
rect 17085 27692 17141 27724
rect 17175 27692 17231 27724
rect 16995 27690 17019 27692
rect 17085 27690 17119 27692
rect 17175 27690 17219 27692
rect 17265 27690 17326 27724
rect 16953 27658 17019 27690
rect 17053 27658 17119 27690
rect 17153 27658 17219 27690
rect 17253 27658 17326 27690
rect 16632 27634 17326 27658
rect 16632 27600 16691 27634
rect 16725 27600 16781 27634
rect 16815 27600 16871 27634
rect 16905 27600 16961 27634
rect 16995 27600 17051 27634
rect 17085 27600 17141 27634
rect 17175 27600 17231 27634
rect 17265 27600 17326 27634
rect 16632 27592 17326 27600
rect 16632 27558 16719 27592
rect 16753 27558 16819 27592
rect 16853 27558 16919 27592
rect 16953 27558 17019 27592
rect 17053 27558 17119 27592
rect 17153 27558 17219 27592
rect 17253 27558 17326 27592
rect 16632 27544 17326 27558
rect 16632 27510 16691 27544
rect 16725 27510 16781 27544
rect 16815 27510 16871 27544
rect 16905 27510 16961 27544
rect 16995 27510 17051 27544
rect 17085 27510 17141 27544
rect 17175 27510 17231 27544
rect 17265 27510 17326 27544
rect 16632 27492 17326 27510
rect 16632 27458 16719 27492
rect 16753 27458 16819 27492
rect 16853 27458 16919 27492
rect 16953 27458 17019 27492
rect 17053 27458 17119 27492
rect 17153 27458 17219 27492
rect 17253 27458 17326 27492
rect 16632 27454 17326 27458
rect 16632 27420 16691 27454
rect 16725 27420 16781 27454
rect 16815 27420 16871 27454
rect 16905 27420 16961 27454
rect 16995 27420 17051 27454
rect 17085 27420 17141 27454
rect 17175 27420 17231 27454
rect 17265 27420 17326 27454
rect 16632 27392 17326 27420
rect 16632 27364 16719 27392
rect 16753 27364 16819 27392
rect 16632 27330 16691 27364
rect 16753 27358 16781 27364
rect 16725 27330 16781 27358
rect 16815 27358 16819 27364
rect 16853 27364 16919 27392
rect 16853 27358 16871 27364
rect 16815 27330 16871 27358
rect 16905 27358 16919 27364
rect 16953 27364 17019 27392
rect 17053 27364 17119 27392
rect 17153 27364 17219 27392
rect 17253 27364 17326 27392
rect 16953 27358 16961 27364
rect 16905 27330 16961 27358
rect 16995 27358 17019 27364
rect 17085 27358 17119 27364
rect 17175 27358 17219 27364
rect 16995 27330 17051 27358
rect 17085 27330 17141 27358
rect 17175 27330 17231 27358
rect 17265 27330 17326 27364
rect 16632 27271 17326 27330
rect 17388 27933 17407 27967
rect 17388 27877 17424 27933
rect 17388 27843 17407 27877
rect 17388 27787 17424 27843
rect 17388 27753 17407 27787
rect 17388 27697 17424 27753
rect 17388 27663 17407 27697
rect 17388 27607 17424 27663
rect 17388 27573 17407 27607
rect 17388 27517 17424 27573
rect 17388 27483 17407 27517
rect 17388 27427 17424 27483
rect 17388 27393 17407 27427
rect 17388 27337 17424 27393
rect 17388 27303 17407 27337
rect 16044 27213 16063 27247
rect 16044 27209 16092 27213
rect 16508 27232 16517 27266
rect 16551 27232 16570 27266
rect 15178 27190 16092 27209
rect 15178 27175 15231 27190
rect 15265 27175 15321 27190
rect 15355 27175 15411 27190
rect 15445 27175 15501 27190
rect 15535 27175 15591 27190
rect 15625 27175 15681 27190
rect 15715 27175 15771 27190
rect 15805 27175 15861 27190
rect 15895 27175 15951 27190
rect 15985 27175 16092 27190
rect 16508 27209 16570 27232
rect 17388 27247 17424 27303
rect 17388 27213 17407 27247
rect 17388 27209 17424 27213
rect 16508 27190 17424 27209
rect 16508 27175 16575 27190
rect 16609 27175 16665 27190
rect 16699 27175 16755 27190
rect 16789 27156 16845 27190
rect 16879 27156 16935 27190
rect 16969 27156 17025 27190
rect 17059 27156 17115 27190
rect 17149 27179 17205 27190
rect 17239 27179 17295 27190
rect 17329 27179 17424 27190
rect 17149 27156 17195 27179
rect 13370 27094 13405 27121
rect 7490 27059 13405 27094
rect 7490 27025 7552 27059
rect 10352 27025 10510 27059
rect 13310 27025 13405 27059
rect 14082 27043 14550 27156
rect 7490 26983 13405 27025
rect 14085 27009 14141 27043
rect 14175 27009 14231 27043
rect 14265 27009 14321 27043
rect 14355 27009 14411 27043
rect 14445 27009 14501 27043
rect 14535 27009 14550 27043
rect 16764 27043 17195 27156
rect 16773 27009 16829 27043
rect 16863 27009 16919 27043
rect 16953 27009 17009 27043
rect 17043 27009 17099 27043
rect 17133 27009 17189 27043
rect 7490 26801 7495 26983
rect 10377 26963 10475 26983
rect 10377 26825 10414 26963
rect 10448 26825 10475 26963
rect 13370 26963 13405 26983
rect 10377 26801 10475 26825
rect 13370 26825 13372 26963
rect 14082 26886 14550 27009
rect 16764 26886 17195 27009
rect 17590 26974 17623 28183
rect 13844 26852 13871 26863
rect 13905 26852 13961 26863
rect 13995 26852 14051 26863
rect 14085 26852 14141 26886
rect 14175 26852 14231 26886
rect 14265 26852 14321 26886
rect 14355 26852 14411 26886
rect 14445 26852 14501 26886
rect 14535 26877 14550 26886
rect 14535 26852 14591 26877
rect 14625 26852 14681 26877
rect 14715 26852 14762 26877
rect 15178 26852 15215 26877
rect 15249 26852 15305 26877
rect 15339 26852 15395 26877
rect 15429 26852 15485 26877
rect 15519 26852 15575 26877
rect 15609 26852 15665 26877
rect 15699 26852 15755 26877
rect 15789 26852 15845 26877
rect 15879 26852 15935 26877
rect 15969 26852 16025 26877
rect 16059 26852 16092 26877
rect 16508 26852 16559 26877
rect 16593 26852 16649 26877
rect 16683 26852 16739 26877
rect 16773 26852 16829 26886
rect 16863 26852 16919 26886
rect 16953 26852 17009 26886
rect 17043 26852 17099 26886
rect 17133 26852 17189 26886
rect 17223 26852 17279 26870
rect 17313 26852 17369 26870
rect 17403 26852 17424 26870
rect 13370 26801 13405 26825
rect 13844 26819 14762 26852
rect 7490 26763 13405 26801
rect 7490 26729 7552 26763
rect 10352 26729 10510 26763
rect 13310 26729 13405 26763
rect 7490 26690 13405 26729
rect 13844 26755 13854 26819
rect 14717 26755 14762 26819
rect 15178 26819 16092 26852
rect 13844 26736 14762 26755
rect 7490 26508 7495 26690
rect 10377 26667 10475 26690
rect 10377 26529 10414 26667
rect 10448 26529 10475 26667
rect 13370 26667 13405 26690
rect 13844 26702 13921 26736
rect 13955 26702 14011 26736
rect 14045 26702 14101 26736
rect 14135 26702 14191 26736
rect 14225 26702 14281 26736
rect 14315 26702 14371 26736
rect 14405 26702 14461 26736
rect 14495 26702 14551 26736
rect 14585 26702 14641 26736
rect 14675 26702 14762 26736
rect 15178 26755 15200 26819
rect 16073 26755 16092 26819
rect 16508 26819 17424 26852
rect 15178 26736 16092 26755
rect 13844 26683 14762 26702
rect 10377 26508 10475 26529
rect 13370 26529 13372 26667
rect 13844 26642 13882 26683
rect 13863 26608 13882 26642
rect 14700 26623 14762 26683
rect 15178 26702 15265 26736
rect 15299 26702 15355 26736
rect 15389 26702 15445 26736
rect 15479 26702 15535 26736
rect 15569 26702 15625 26736
rect 15659 26702 15715 26736
rect 15749 26702 15805 26736
rect 15839 26702 15895 26736
rect 15929 26702 15985 26736
rect 16019 26702 16092 26736
rect 16508 26755 16533 26819
rect 17416 26755 17424 26819
rect 16508 26736 17424 26755
rect 15178 26683 16092 26702
rect 15178 26642 15226 26683
rect 13844 26552 13882 26608
rect 13370 26508 13405 26529
rect 7490 26467 13405 26508
rect 13863 26518 13882 26552
rect 7490 26433 7552 26467
rect 10352 26433 10510 26467
rect 13310 26433 13405 26467
rect 13844 26462 13882 26518
rect 7490 26397 13405 26433
rect 13863 26428 13882 26462
rect 7490 26208 7495 26397
rect 10377 26371 10475 26397
rect 10377 26233 10414 26371
rect 10448 26233 10475 26371
rect 13370 26371 13405 26397
rect 13844 26372 13882 26428
rect 10377 26208 10475 26233
rect 13370 26233 13372 26371
rect 13863 26338 13882 26372
rect 13844 26282 13882 26338
rect 13370 26208 13405 26233
rect 13863 26248 13882 26282
rect 7490 26171 13405 26208
rect 13844 26192 13882 26248
rect 7490 26137 7552 26171
rect 10352 26137 10510 26171
rect 13310 26137 13405 26171
rect 13863 26158 13882 26192
rect 7490 26097 13405 26137
rect 13844 26102 13882 26158
rect 7490 25901 7495 26097
rect 10377 26075 10475 26097
rect 10377 25937 10414 26075
rect 10448 25937 10475 26075
rect 13370 26075 13405 26097
rect 10377 25901 10475 25937
rect 13370 25937 13372 26075
rect 13863 26068 13882 26102
rect 13844 26012 13882 26068
rect 13863 25978 13882 26012
rect 13370 25901 13405 25937
rect 13844 25922 13882 25978
rect 13944 26560 14638 26621
rect 13944 26526 14003 26560
rect 14037 26548 14093 26560
rect 14065 26526 14093 26548
rect 14127 26548 14183 26560
rect 14127 26526 14131 26548
rect 13944 26514 14031 26526
rect 14065 26514 14131 26526
rect 14165 26526 14183 26548
rect 14217 26548 14273 26560
rect 14217 26526 14231 26548
rect 14165 26514 14231 26526
rect 14265 26526 14273 26548
rect 14307 26548 14363 26560
rect 14397 26548 14453 26560
rect 14487 26548 14543 26560
rect 14307 26526 14331 26548
rect 14397 26526 14431 26548
rect 14487 26526 14531 26548
rect 14577 26526 14638 26560
rect 14265 26514 14331 26526
rect 14365 26514 14431 26526
rect 14465 26514 14531 26526
rect 14565 26514 14638 26526
rect 13944 26470 14638 26514
rect 13944 26436 14003 26470
rect 14037 26448 14093 26470
rect 14065 26436 14093 26448
rect 14127 26448 14183 26470
rect 14127 26436 14131 26448
rect 13944 26414 14031 26436
rect 14065 26414 14131 26436
rect 14165 26436 14183 26448
rect 14217 26448 14273 26470
rect 14217 26436 14231 26448
rect 14165 26414 14231 26436
rect 14265 26436 14273 26448
rect 14307 26448 14363 26470
rect 14397 26448 14453 26470
rect 14487 26448 14543 26470
rect 14307 26436 14331 26448
rect 14397 26436 14431 26448
rect 14487 26436 14531 26448
rect 14577 26436 14638 26470
rect 14265 26414 14331 26436
rect 14365 26414 14431 26436
rect 14465 26414 14531 26436
rect 14565 26414 14638 26436
rect 13944 26380 14638 26414
rect 13944 26346 14003 26380
rect 14037 26348 14093 26380
rect 14065 26346 14093 26348
rect 14127 26348 14183 26380
rect 14127 26346 14131 26348
rect 13944 26314 14031 26346
rect 14065 26314 14131 26346
rect 14165 26346 14183 26348
rect 14217 26348 14273 26380
rect 14217 26346 14231 26348
rect 14165 26314 14231 26346
rect 14265 26346 14273 26348
rect 14307 26348 14363 26380
rect 14397 26348 14453 26380
rect 14487 26348 14543 26380
rect 14307 26346 14331 26348
rect 14397 26346 14431 26348
rect 14487 26346 14531 26348
rect 14577 26346 14638 26380
rect 14265 26314 14331 26346
rect 14365 26314 14431 26346
rect 14465 26314 14531 26346
rect 14565 26314 14638 26346
rect 13944 26290 14638 26314
rect 13944 26256 14003 26290
rect 14037 26256 14093 26290
rect 14127 26256 14183 26290
rect 14217 26256 14273 26290
rect 14307 26256 14363 26290
rect 14397 26256 14453 26290
rect 14487 26256 14543 26290
rect 14577 26256 14638 26290
rect 13944 26248 14638 26256
rect 13944 26214 14031 26248
rect 14065 26214 14131 26248
rect 14165 26214 14231 26248
rect 14265 26214 14331 26248
rect 14365 26214 14431 26248
rect 14465 26214 14531 26248
rect 14565 26214 14638 26248
rect 13944 26200 14638 26214
rect 13944 26166 14003 26200
rect 14037 26166 14093 26200
rect 14127 26166 14183 26200
rect 14217 26166 14273 26200
rect 14307 26166 14363 26200
rect 14397 26166 14453 26200
rect 14487 26166 14543 26200
rect 14577 26166 14638 26200
rect 13944 26148 14638 26166
rect 13944 26114 14031 26148
rect 14065 26114 14131 26148
rect 14165 26114 14231 26148
rect 14265 26114 14331 26148
rect 14365 26114 14431 26148
rect 14465 26114 14531 26148
rect 14565 26114 14638 26148
rect 13944 26110 14638 26114
rect 13944 26076 14003 26110
rect 14037 26076 14093 26110
rect 14127 26076 14183 26110
rect 14217 26076 14273 26110
rect 14307 26076 14363 26110
rect 14397 26076 14453 26110
rect 14487 26076 14543 26110
rect 14577 26076 14638 26110
rect 13944 26048 14638 26076
rect 13944 26020 14031 26048
rect 14065 26020 14131 26048
rect 13944 25986 14003 26020
rect 14065 26014 14093 26020
rect 14037 25986 14093 26014
rect 14127 26014 14131 26020
rect 14165 26020 14231 26048
rect 14165 26014 14183 26020
rect 14127 25986 14183 26014
rect 14217 26014 14231 26020
rect 14265 26020 14331 26048
rect 14365 26020 14431 26048
rect 14465 26020 14531 26048
rect 14565 26020 14638 26048
rect 14265 26014 14273 26020
rect 14217 25986 14273 26014
rect 14307 26014 14331 26020
rect 14397 26014 14431 26020
rect 14487 26014 14531 26020
rect 14307 25986 14363 26014
rect 14397 25986 14453 26014
rect 14487 25986 14543 26014
rect 14577 25986 14638 26020
rect 13944 25927 14638 25986
rect 14700 26589 14719 26623
rect 14753 26589 14762 26623
rect 14700 26533 14762 26589
rect 15207 26608 15226 26642
rect 16044 26623 16092 26683
rect 16508 26702 16609 26736
rect 16643 26702 16699 26736
rect 16733 26702 16789 26736
rect 16823 26702 16879 26736
rect 16913 26702 16969 26736
rect 17003 26702 17059 26736
rect 17093 26702 17149 26736
rect 17183 26702 17239 26736
rect 17273 26702 17329 26736
rect 17363 26702 17424 26736
rect 16508 26683 17424 26702
rect 16508 26642 16570 26683
rect 15178 26552 15226 26608
rect 14700 26499 14719 26533
rect 14753 26499 14762 26533
rect 14700 26443 14762 26499
rect 15207 26518 15226 26552
rect 15178 26462 15226 26518
rect 14700 26409 14719 26443
rect 14753 26409 14762 26443
rect 14700 26353 14762 26409
rect 15207 26428 15226 26462
rect 15178 26372 15226 26428
rect 14700 26319 14719 26353
rect 14753 26319 14762 26353
rect 14700 26263 14762 26319
rect 15207 26338 15226 26372
rect 15178 26282 15226 26338
rect 14700 26229 14719 26263
rect 14753 26229 14762 26263
rect 14700 26173 14762 26229
rect 15207 26248 15226 26282
rect 15178 26192 15226 26248
rect 14700 26139 14719 26173
rect 14753 26139 14762 26173
rect 14700 26083 14762 26139
rect 15207 26158 15226 26192
rect 15178 26102 15226 26158
rect 14700 26049 14719 26083
rect 14753 26049 14762 26083
rect 14700 25993 14762 26049
rect 15207 26068 15226 26102
rect 15178 26012 15226 26068
rect 14700 25959 14719 25993
rect 14753 25959 14762 25993
rect 7490 25875 13405 25901
rect 7490 25841 7552 25875
rect 10352 25841 10510 25875
rect 13310 25841 13405 25875
rect 13863 25888 13882 25922
rect 7490 25790 13405 25841
rect 13844 25865 13882 25888
rect 14700 25903 14762 25959
rect 15207 25978 15226 26012
rect 15178 25922 15226 25978
rect 15288 26560 15982 26621
rect 15288 26526 15347 26560
rect 15381 26548 15437 26560
rect 15409 26526 15437 26548
rect 15471 26548 15527 26560
rect 15471 26526 15475 26548
rect 15288 26514 15375 26526
rect 15409 26514 15475 26526
rect 15509 26526 15527 26548
rect 15561 26548 15617 26560
rect 15561 26526 15575 26548
rect 15509 26514 15575 26526
rect 15609 26526 15617 26548
rect 15651 26548 15707 26560
rect 15741 26548 15797 26560
rect 15831 26548 15887 26560
rect 15651 26526 15675 26548
rect 15741 26526 15775 26548
rect 15831 26526 15875 26548
rect 15921 26526 15982 26560
rect 15609 26514 15675 26526
rect 15709 26514 15775 26526
rect 15809 26514 15875 26526
rect 15909 26514 15982 26526
rect 15288 26470 15982 26514
rect 15288 26436 15347 26470
rect 15381 26448 15437 26470
rect 15409 26436 15437 26448
rect 15471 26448 15527 26470
rect 15471 26436 15475 26448
rect 15288 26414 15375 26436
rect 15409 26414 15475 26436
rect 15509 26436 15527 26448
rect 15561 26448 15617 26470
rect 15561 26436 15575 26448
rect 15509 26414 15575 26436
rect 15609 26436 15617 26448
rect 15651 26448 15707 26470
rect 15741 26448 15797 26470
rect 15831 26448 15887 26470
rect 15651 26436 15675 26448
rect 15741 26436 15775 26448
rect 15831 26436 15875 26448
rect 15921 26436 15982 26470
rect 15609 26414 15675 26436
rect 15709 26414 15775 26436
rect 15809 26414 15875 26436
rect 15909 26414 15982 26436
rect 15288 26380 15982 26414
rect 15288 26346 15347 26380
rect 15381 26348 15437 26380
rect 15409 26346 15437 26348
rect 15471 26348 15527 26380
rect 15471 26346 15475 26348
rect 15288 26314 15375 26346
rect 15409 26314 15475 26346
rect 15509 26346 15527 26348
rect 15561 26348 15617 26380
rect 15561 26346 15575 26348
rect 15509 26314 15575 26346
rect 15609 26346 15617 26348
rect 15651 26348 15707 26380
rect 15741 26348 15797 26380
rect 15831 26348 15887 26380
rect 15651 26346 15675 26348
rect 15741 26346 15775 26348
rect 15831 26346 15875 26348
rect 15921 26346 15982 26380
rect 15609 26314 15675 26346
rect 15709 26314 15775 26346
rect 15809 26314 15875 26346
rect 15909 26314 15982 26346
rect 15288 26290 15982 26314
rect 15288 26256 15347 26290
rect 15381 26256 15437 26290
rect 15471 26256 15527 26290
rect 15561 26256 15617 26290
rect 15651 26256 15707 26290
rect 15741 26256 15797 26290
rect 15831 26256 15887 26290
rect 15921 26256 15982 26290
rect 15288 26248 15982 26256
rect 15288 26214 15375 26248
rect 15409 26214 15475 26248
rect 15509 26214 15575 26248
rect 15609 26214 15675 26248
rect 15709 26214 15775 26248
rect 15809 26214 15875 26248
rect 15909 26214 15982 26248
rect 15288 26200 15982 26214
rect 15288 26166 15347 26200
rect 15381 26166 15437 26200
rect 15471 26166 15527 26200
rect 15561 26166 15617 26200
rect 15651 26166 15707 26200
rect 15741 26166 15797 26200
rect 15831 26166 15887 26200
rect 15921 26166 15982 26200
rect 15288 26148 15982 26166
rect 15288 26114 15375 26148
rect 15409 26114 15475 26148
rect 15509 26114 15575 26148
rect 15609 26114 15675 26148
rect 15709 26114 15775 26148
rect 15809 26114 15875 26148
rect 15909 26114 15982 26148
rect 15288 26110 15982 26114
rect 15288 26076 15347 26110
rect 15381 26076 15437 26110
rect 15471 26076 15527 26110
rect 15561 26076 15617 26110
rect 15651 26076 15707 26110
rect 15741 26076 15797 26110
rect 15831 26076 15887 26110
rect 15921 26076 15982 26110
rect 15288 26048 15982 26076
rect 15288 26020 15375 26048
rect 15409 26020 15475 26048
rect 15288 25986 15347 26020
rect 15409 26014 15437 26020
rect 15381 25986 15437 26014
rect 15471 26014 15475 26020
rect 15509 26020 15575 26048
rect 15509 26014 15527 26020
rect 15471 25986 15527 26014
rect 15561 26014 15575 26020
rect 15609 26020 15675 26048
rect 15709 26020 15775 26048
rect 15809 26020 15875 26048
rect 15909 26020 15982 26048
rect 15609 26014 15617 26020
rect 15561 25986 15617 26014
rect 15651 26014 15675 26020
rect 15741 26014 15775 26020
rect 15831 26014 15875 26020
rect 15651 25986 15707 26014
rect 15741 25986 15797 26014
rect 15831 25986 15887 26014
rect 15921 25986 15982 26020
rect 15288 25927 15982 25986
rect 16044 26589 16063 26623
rect 16044 26533 16092 26589
rect 16508 26608 16517 26642
rect 16551 26608 16570 26642
rect 17388 26623 17424 26683
rect 16508 26552 16570 26608
rect 16044 26499 16063 26533
rect 16044 26443 16092 26499
rect 16508 26518 16517 26552
rect 16551 26518 16570 26552
rect 16508 26462 16570 26518
rect 16044 26409 16063 26443
rect 16044 26353 16092 26409
rect 16508 26428 16517 26462
rect 16551 26428 16570 26462
rect 16508 26372 16570 26428
rect 16044 26319 16063 26353
rect 16044 26263 16092 26319
rect 16508 26338 16517 26372
rect 16551 26338 16570 26372
rect 16508 26282 16570 26338
rect 16044 26229 16063 26263
rect 16044 26173 16092 26229
rect 16508 26248 16517 26282
rect 16551 26248 16570 26282
rect 16508 26192 16570 26248
rect 16044 26139 16063 26173
rect 16044 26083 16092 26139
rect 16508 26158 16517 26192
rect 16551 26158 16570 26192
rect 16508 26102 16570 26158
rect 16044 26049 16063 26083
rect 16044 25993 16092 26049
rect 16508 26068 16517 26102
rect 16551 26068 16570 26102
rect 16508 26012 16570 26068
rect 16044 25959 16063 25993
rect 14700 25869 14719 25903
rect 14753 25869 14762 25903
rect 14700 25865 14762 25869
rect 15207 25888 15226 25922
rect 13844 25846 14762 25865
rect 13844 25826 13887 25846
rect 13921 25826 13977 25846
rect 14011 25826 14067 25846
rect 14101 25812 14157 25846
rect 14191 25812 14247 25846
rect 14281 25812 14337 25846
rect 14371 25812 14427 25846
rect 14461 25812 14517 25846
rect 14551 25826 14607 25846
rect 14641 25826 14762 25846
rect 15178 25865 15226 25888
rect 16044 25903 16092 25959
rect 16508 25978 16517 26012
rect 16551 25978 16570 26012
rect 16508 25922 16570 25978
rect 16632 26560 17326 26621
rect 16632 26526 16691 26560
rect 16725 26548 16781 26560
rect 16753 26526 16781 26548
rect 16815 26548 16871 26560
rect 16815 26526 16819 26548
rect 16632 26514 16719 26526
rect 16753 26514 16819 26526
rect 16853 26526 16871 26548
rect 16905 26548 16961 26560
rect 16905 26526 16919 26548
rect 16853 26514 16919 26526
rect 16953 26526 16961 26548
rect 16995 26548 17051 26560
rect 17085 26548 17141 26560
rect 17175 26548 17231 26560
rect 16995 26526 17019 26548
rect 17085 26526 17119 26548
rect 17175 26526 17219 26548
rect 17265 26526 17326 26560
rect 16953 26514 17019 26526
rect 17053 26514 17119 26526
rect 17153 26514 17219 26526
rect 17253 26514 17326 26526
rect 16632 26470 17326 26514
rect 16632 26436 16691 26470
rect 16725 26448 16781 26470
rect 16753 26436 16781 26448
rect 16815 26448 16871 26470
rect 16815 26436 16819 26448
rect 16632 26414 16719 26436
rect 16753 26414 16819 26436
rect 16853 26436 16871 26448
rect 16905 26448 16961 26470
rect 16905 26436 16919 26448
rect 16853 26414 16919 26436
rect 16953 26436 16961 26448
rect 16995 26448 17051 26470
rect 17085 26448 17141 26470
rect 17175 26448 17231 26470
rect 16995 26436 17019 26448
rect 17085 26436 17119 26448
rect 17175 26436 17219 26448
rect 17265 26436 17326 26470
rect 16953 26414 17019 26436
rect 17053 26414 17119 26436
rect 17153 26414 17219 26436
rect 17253 26414 17326 26436
rect 16632 26380 17326 26414
rect 16632 26346 16691 26380
rect 16725 26348 16781 26380
rect 16753 26346 16781 26348
rect 16815 26348 16871 26380
rect 16815 26346 16819 26348
rect 16632 26314 16719 26346
rect 16753 26314 16819 26346
rect 16853 26346 16871 26348
rect 16905 26348 16961 26380
rect 16905 26346 16919 26348
rect 16853 26314 16919 26346
rect 16953 26346 16961 26348
rect 16995 26348 17051 26380
rect 17085 26348 17141 26380
rect 17175 26348 17231 26380
rect 16995 26346 17019 26348
rect 17085 26346 17119 26348
rect 17175 26346 17219 26348
rect 17265 26346 17326 26380
rect 16953 26314 17019 26346
rect 17053 26314 17119 26346
rect 17153 26314 17219 26346
rect 17253 26314 17326 26346
rect 16632 26290 17326 26314
rect 16632 26256 16691 26290
rect 16725 26256 16781 26290
rect 16815 26256 16871 26290
rect 16905 26256 16961 26290
rect 16995 26256 17051 26290
rect 17085 26256 17141 26290
rect 17175 26256 17231 26290
rect 17265 26256 17326 26290
rect 16632 26248 17326 26256
rect 16632 26214 16719 26248
rect 16753 26214 16819 26248
rect 16853 26214 16919 26248
rect 16953 26214 17019 26248
rect 17053 26214 17119 26248
rect 17153 26214 17219 26248
rect 17253 26214 17326 26248
rect 16632 26200 17326 26214
rect 16632 26166 16691 26200
rect 16725 26166 16781 26200
rect 16815 26166 16871 26200
rect 16905 26166 16961 26200
rect 16995 26166 17051 26200
rect 17085 26166 17141 26200
rect 17175 26166 17231 26200
rect 17265 26166 17326 26200
rect 16632 26148 17326 26166
rect 16632 26114 16719 26148
rect 16753 26114 16819 26148
rect 16853 26114 16919 26148
rect 16953 26114 17019 26148
rect 17053 26114 17119 26148
rect 17153 26114 17219 26148
rect 17253 26114 17326 26148
rect 16632 26110 17326 26114
rect 16632 26076 16691 26110
rect 16725 26076 16781 26110
rect 16815 26076 16871 26110
rect 16905 26076 16961 26110
rect 16995 26076 17051 26110
rect 17085 26076 17141 26110
rect 17175 26076 17231 26110
rect 17265 26076 17326 26110
rect 16632 26048 17326 26076
rect 16632 26020 16719 26048
rect 16753 26020 16819 26048
rect 16632 25986 16691 26020
rect 16753 26014 16781 26020
rect 16725 25986 16781 26014
rect 16815 26014 16819 26020
rect 16853 26020 16919 26048
rect 16853 26014 16871 26020
rect 16815 25986 16871 26014
rect 16905 26014 16919 26020
rect 16953 26020 17019 26048
rect 17053 26020 17119 26048
rect 17153 26020 17219 26048
rect 17253 26020 17326 26048
rect 16953 26014 16961 26020
rect 16905 25986 16961 26014
rect 16995 26014 17019 26020
rect 17085 26014 17119 26020
rect 17175 26014 17219 26020
rect 16995 25986 17051 26014
rect 17085 25986 17141 26014
rect 17175 25986 17231 26014
rect 17265 25986 17326 26020
rect 16632 25927 17326 25986
rect 17388 26589 17407 26623
rect 17388 26533 17424 26589
rect 17388 26499 17407 26533
rect 17388 26443 17424 26499
rect 17388 26409 17407 26443
rect 17388 26353 17424 26409
rect 17388 26319 17407 26353
rect 17388 26263 17424 26319
rect 17388 26229 17407 26263
rect 17388 26173 17424 26229
rect 17388 26139 17407 26173
rect 17388 26083 17424 26139
rect 17388 26049 17407 26083
rect 17388 25993 17424 26049
rect 17388 25959 17407 25993
rect 16044 25869 16063 25903
rect 16044 25865 16092 25869
rect 16508 25888 16517 25922
rect 16551 25888 16570 25922
rect 15178 25846 16092 25865
rect 15178 25826 15231 25846
rect 15265 25826 15321 25846
rect 15355 25826 15411 25846
rect 15445 25826 15501 25846
rect 15535 25826 15591 25846
rect 15625 25826 15681 25846
rect 15715 25826 15771 25846
rect 15805 25826 15861 25846
rect 15895 25826 15951 25846
rect 15985 25826 16092 25846
rect 16508 25865 16570 25888
rect 17388 25903 17424 25959
rect 17388 25869 17407 25903
rect 17388 25865 17424 25869
rect 16508 25846 17424 25865
rect 16508 25826 16575 25846
rect 16609 25826 16665 25846
rect 16699 25826 16755 25846
rect 14551 25812 14581 25826
rect 16753 25812 16755 25826
rect 16789 25812 16845 25846
rect 16879 25812 16935 25846
rect 16969 25812 17025 25846
rect 17059 25812 17115 25846
rect 17149 25812 17205 25846
rect 17239 25845 17295 25846
rect 17329 25845 17424 25846
rect 7490 25615 7495 25790
rect 10377 25779 10475 25790
rect 10377 25641 10414 25779
rect 10448 25641 10475 25779
rect 13370 25779 13405 25790
rect 10377 25615 10475 25641
rect 13370 25641 13372 25779
rect 14082 25699 14581 25812
rect 14085 25665 14141 25699
rect 14175 25665 14231 25699
rect 14265 25665 14321 25699
rect 14355 25665 14411 25699
rect 14445 25665 14501 25699
rect 14535 25665 14581 25699
rect 16753 25699 17210 25812
rect 16773 25665 16829 25699
rect 16863 25665 16919 25699
rect 16953 25665 17009 25699
rect 17043 25665 17099 25699
rect 17133 25665 17189 25699
rect 13370 25615 13405 25641
rect 7490 25579 13405 25615
rect 7490 25545 7552 25579
rect 10352 25545 10510 25579
rect 13310 25545 13405 25579
rect 7490 25504 13405 25545
rect 14082 25542 14581 25665
rect 16753 25542 17210 25665
rect 17590 25630 17623 26918
rect 13844 25508 13871 25517
rect 13905 25508 13961 25517
rect 13995 25508 14051 25517
rect 14085 25508 14141 25542
rect 14175 25508 14231 25542
rect 14265 25508 14321 25542
rect 14355 25508 14411 25542
rect 14445 25508 14501 25542
rect 14535 25520 14581 25542
rect 14535 25508 14591 25520
rect 14625 25508 14681 25520
rect 14715 25508 14762 25520
rect 15178 25508 15215 25520
rect 15249 25508 15305 25520
rect 15339 25508 15395 25520
rect 15429 25508 15485 25520
rect 15519 25508 15575 25520
rect 15609 25508 15665 25520
rect 15699 25508 15755 25520
rect 15789 25508 15845 25520
rect 15879 25508 15935 25520
rect 15969 25508 16025 25520
rect 16059 25508 16092 25520
rect 16508 25508 16559 25520
rect 16593 25508 16649 25520
rect 16683 25508 16739 25520
rect 16773 25508 16829 25542
rect 16863 25508 16919 25542
rect 16953 25508 17009 25542
rect 17043 25508 17099 25542
rect 17133 25508 17189 25542
rect 7490 25322 7495 25504
rect 10377 25483 10475 25504
rect 10377 25345 10414 25483
rect 10448 25345 10475 25483
rect 13370 25483 13405 25504
rect 10377 25322 10475 25345
rect 13370 25345 13372 25483
rect 13844 25392 14762 25508
rect 13370 25322 13405 25345
rect 13844 25358 13921 25392
rect 13955 25358 14011 25392
rect 14045 25358 14101 25392
rect 14135 25358 14191 25392
rect 14225 25358 14281 25392
rect 14315 25358 14371 25392
rect 14405 25358 14461 25392
rect 14495 25358 14551 25392
rect 14585 25358 14641 25392
rect 14675 25358 14762 25392
rect 15178 25392 16092 25508
rect 16508 25501 17210 25508
rect 13844 25339 14762 25358
rect 7490 25283 13405 25322
rect 13844 25298 13882 25339
rect 7490 25249 7552 25283
rect 10352 25249 10510 25283
rect 13310 25249 13405 25283
rect 7490 25211 13405 25249
rect 13863 25264 13882 25298
rect 14700 25279 14762 25339
rect 15178 25358 15265 25392
rect 15299 25358 15355 25392
rect 15389 25358 15445 25392
rect 15479 25358 15535 25392
rect 15569 25358 15625 25392
rect 15659 25358 15715 25392
rect 15749 25358 15805 25392
rect 15839 25358 15895 25392
rect 15929 25358 15985 25392
rect 16019 25358 16092 25392
rect 16508 25392 17424 25501
rect 15178 25339 16092 25358
rect 15178 25298 15226 25339
rect 7490 25015 7495 25211
rect 10377 25187 10475 25211
rect 10377 25049 10414 25187
rect 10448 25049 10475 25187
rect 13370 25187 13405 25211
rect 13844 25208 13882 25264
rect 10377 25015 10475 25049
rect 13370 25049 13372 25187
rect 13863 25174 13882 25208
rect 13844 25118 13882 25174
rect 13863 25084 13882 25118
rect 13370 25015 13405 25049
rect 13844 25028 13882 25084
rect 7490 24987 13405 25015
rect 7490 24953 7552 24987
rect 10352 24953 10510 24987
rect 13310 24953 13405 24987
rect 13863 24994 13882 25028
rect 7490 24904 13405 24953
rect 13844 24938 13882 24994
rect 5742 24621 7371 24690
rect 5981 24614 7371 24621
rect 7490 24701 7495 24904
rect 10377 24891 10475 24904
rect 10377 24753 10414 24891
rect 10448 24753 10475 24891
rect 13370 24891 13405 24904
rect 10377 24701 10475 24753
rect 13370 24753 13372 24891
rect 13863 24904 13882 24938
rect 13844 24848 13882 24904
rect 13863 24814 13882 24848
rect 13844 24758 13882 24814
rect 13370 24701 13405 24753
rect 13863 24724 13882 24758
rect 7490 24691 13405 24701
rect 7490 24657 7552 24691
rect 10352 24657 10510 24691
rect 13310 24657 13405 24691
rect 13844 24668 13882 24724
rect 7490 24614 13405 24657
rect 13863 24634 13882 24668
rect 11232 24602 13405 24614
rect 13844 24578 13882 24634
rect 13944 25216 14638 25277
rect 13944 25182 14003 25216
rect 14037 25204 14093 25216
rect 14065 25182 14093 25204
rect 14127 25204 14183 25216
rect 14127 25182 14131 25204
rect 13944 25170 14031 25182
rect 14065 25170 14131 25182
rect 14165 25182 14183 25204
rect 14217 25204 14273 25216
rect 14217 25182 14231 25204
rect 14165 25170 14231 25182
rect 14265 25182 14273 25204
rect 14307 25204 14363 25216
rect 14397 25204 14453 25216
rect 14487 25204 14543 25216
rect 14307 25182 14331 25204
rect 14397 25182 14431 25204
rect 14487 25182 14531 25204
rect 14577 25182 14638 25216
rect 14265 25170 14331 25182
rect 14365 25170 14431 25182
rect 14465 25170 14531 25182
rect 14565 25170 14638 25182
rect 13944 25126 14638 25170
rect 13944 25092 14003 25126
rect 14037 25104 14093 25126
rect 14065 25092 14093 25104
rect 14127 25104 14183 25126
rect 14127 25092 14131 25104
rect 13944 25070 14031 25092
rect 14065 25070 14131 25092
rect 14165 25092 14183 25104
rect 14217 25104 14273 25126
rect 14217 25092 14231 25104
rect 14165 25070 14231 25092
rect 14265 25092 14273 25104
rect 14307 25104 14363 25126
rect 14397 25104 14453 25126
rect 14487 25104 14543 25126
rect 14307 25092 14331 25104
rect 14397 25092 14431 25104
rect 14487 25092 14531 25104
rect 14577 25092 14638 25126
rect 14265 25070 14331 25092
rect 14365 25070 14431 25092
rect 14465 25070 14531 25092
rect 14565 25070 14638 25092
rect 13944 25036 14638 25070
rect 13944 25002 14003 25036
rect 14037 25004 14093 25036
rect 14065 25002 14093 25004
rect 14127 25004 14183 25036
rect 14127 25002 14131 25004
rect 13944 24970 14031 25002
rect 14065 24970 14131 25002
rect 14165 25002 14183 25004
rect 14217 25004 14273 25036
rect 14217 25002 14231 25004
rect 14165 24970 14231 25002
rect 14265 25002 14273 25004
rect 14307 25004 14363 25036
rect 14397 25004 14453 25036
rect 14487 25004 14543 25036
rect 14307 25002 14331 25004
rect 14397 25002 14431 25004
rect 14487 25002 14531 25004
rect 14577 25002 14638 25036
rect 14265 24970 14331 25002
rect 14365 24970 14431 25002
rect 14465 24970 14531 25002
rect 14565 24970 14638 25002
rect 13944 24946 14638 24970
rect 13944 24912 14003 24946
rect 14037 24912 14093 24946
rect 14127 24912 14183 24946
rect 14217 24912 14273 24946
rect 14307 24912 14363 24946
rect 14397 24912 14453 24946
rect 14487 24912 14543 24946
rect 14577 24912 14638 24946
rect 13944 24904 14638 24912
rect 13944 24870 14031 24904
rect 14065 24870 14131 24904
rect 14165 24870 14231 24904
rect 14265 24870 14331 24904
rect 14365 24870 14431 24904
rect 14465 24870 14531 24904
rect 14565 24870 14638 24904
rect 13944 24856 14638 24870
rect 13944 24822 14003 24856
rect 14037 24822 14093 24856
rect 14127 24822 14183 24856
rect 14217 24822 14273 24856
rect 14307 24822 14363 24856
rect 14397 24822 14453 24856
rect 14487 24822 14543 24856
rect 14577 24822 14638 24856
rect 13944 24804 14638 24822
rect 13944 24770 14031 24804
rect 14065 24770 14131 24804
rect 14165 24770 14231 24804
rect 14265 24770 14331 24804
rect 14365 24770 14431 24804
rect 14465 24770 14531 24804
rect 14565 24770 14638 24804
rect 13944 24766 14638 24770
rect 13944 24732 14003 24766
rect 14037 24732 14093 24766
rect 14127 24732 14183 24766
rect 14217 24732 14273 24766
rect 14307 24732 14363 24766
rect 14397 24732 14453 24766
rect 14487 24732 14543 24766
rect 14577 24732 14638 24766
rect 13944 24704 14638 24732
rect 13944 24676 14031 24704
rect 14065 24676 14131 24704
rect 13944 24642 14003 24676
rect 14065 24670 14093 24676
rect 14037 24642 14093 24670
rect 14127 24670 14131 24676
rect 14165 24676 14231 24704
rect 14165 24670 14183 24676
rect 14127 24642 14183 24670
rect 14217 24670 14231 24676
rect 14265 24676 14331 24704
rect 14365 24676 14431 24704
rect 14465 24676 14531 24704
rect 14565 24676 14638 24704
rect 14265 24670 14273 24676
rect 14217 24642 14273 24670
rect 14307 24670 14331 24676
rect 14397 24670 14431 24676
rect 14487 24670 14531 24676
rect 14307 24642 14363 24670
rect 14397 24642 14453 24670
rect 14487 24642 14543 24670
rect 14577 24642 14638 24676
rect 13944 24583 14638 24642
rect 14700 25245 14719 25279
rect 14753 25245 14762 25279
rect 14700 25189 14762 25245
rect 15207 25264 15226 25298
rect 16044 25279 16092 25339
rect 16508 25358 16609 25392
rect 16643 25358 16699 25392
rect 16733 25358 16789 25392
rect 16823 25358 16879 25392
rect 16913 25358 16969 25392
rect 17003 25358 17059 25392
rect 17093 25358 17149 25392
rect 17183 25358 17239 25392
rect 17273 25358 17329 25392
rect 17363 25358 17424 25392
rect 16508 25339 17424 25358
rect 16508 25298 16570 25339
rect 15178 25208 15226 25264
rect 14700 25155 14719 25189
rect 14753 25155 14762 25189
rect 14700 25105 14762 25155
rect 15207 25174 15226 25208
rect 15178 25118 15226 25174
rect 14700 25099 15173 25105
rect 14700 25065 14719 25099
rect 14753 25098 15173 25099
rect 14753 25065 14867 25098
rect 14700 25064 14867 25065
rect 14901 25064 15024 25098
rect 15058 25084 15173 25098
rect 15207 25084 15226 25118
rect 15058 25064 15226 25084
rect 14700 25028 15226 25064
rect 14700 25009 15173 25028
rect 14700 24975 14719 25009
rect 14753 25008 15173 25009
rect 14753 24975 14867 25008
rect 14700 24974 14867 24975
rect 14901 24974 15024 25008
rect 15058 24994 15173 25008
rect 15207 24994 15226 25028
rect 15058 24974 15226 24994
rect 14700 24938 15226 24974
rect 14700 24919 15173 24938
rect 14700 24885 14719 24919
rect 14753 24918 15173 24919
rect 14753 24885 14867 24918
rect 14700 24884 14867 24885
rect 14901 24884 15024 24918
rect 15058 24904 15173 24918
rect 15207 24904 15226 24938
rect 15058 24884 15226 24904
rect 14700 24848 15226 24884
rect 14700 24829 15173 24848
rect 14700 24795 14719 24829
rect 14753 24828 15173 24829
rect 14753 24795 14867 24828
rect 14700 24794 14867 24795
rect 14901 24794 15024 24828
rect 15058 24814 15173 24828
rect 15207 24814 15226 24848
rect 15058 24794 15226 24814
rect 14700 24758 15226 24794
rect 14700 24739 15173 24758
rect 14700 24705 14719 24739
rect 14753 24738 15173 24739
rect 14753 24716 14867 24738
rect 14901 24716 15024 24738
rect 15058 24724 15173 24738
rect 15207 24724 15226 24758
rect 15058 24716 15226 24724
rect 14700 24649 14743 24705
rect 15185 24668 15226 24716
rect 14700 24615 14719 24649
rect 13863 24544 13882 24578
rect 13844 24521 13882 24544
rect 14700 24559 14743 24615
rect 15207 24634 15226 24668
rect 15185 24578 15226 24634
rect 15288 25216 15982 25277
rect 15288 25182 15347 25216
rect 15381 25204 15437 25216
rect 15409 25182 15437 25204
rect 15471 25204 15527 25216
rect 15471 25182 15475 25204
rect 15288 25170 15375 25182
rect 15409 25170 15475 25182
rect 15509 25182 15527 25204
rect 15561 25204 15617 25216
rect 15561 25182 15575 25204
rect 15509 25170 15575 25182
rect 15609 25182 15617 25204
rect 15651 25204 15707 25216
rect 15741 25204 15797 25216
rect 15831 25204 15887 25216
rect 15651 25182 15675 25204
rect 15741 25182 15775 25204
rect 15831 25182 15875 25204
rect 15921 25182 15982 25216
rect 15609 25170 15675 25182
rect 15709 25170 15775 25182
rect 15809 25170 15875 25182
rect 15909 25170 15982 25182
rect 15288 25126 15982 25170
rect 15288 25092 15347 25126
rect 15381 25104 15437 25126
rect 15409 25092 15437 25104
rect 15471 25104 15527 25126
rect 15471 25092 15475 25104
rect 15288 25070 15375 25092
rect 15409 25070 15475 25092
rect 15509 25092 15527 25104
rect 15561 25104 15617 25126
rect 15561 25092 15575 25104
rect 15509 25070 15575 25092
rect 15609 25092 15617 25104
rect 15651 25104 15707 25126
rect 15741 25104 15797 25126
rect 15831 25104 15887 25126
rect 15651 25092 15675 25104
rect 15741 25092 15775 25104
rect 15831 25092 15875 25104
rect 15921 25092 15982 25126
rect 15609 25070 15675 25092
rect 15709 25070 15775 25092
rect 15809 25070 15875 25092
rect 15909 25070 15982 25092
rect 15288 25036 15982 25070
rect 15288 25002 15347 25036
rect 15381 25004 15437 25036
rect 15409 25002 15437 25004
rect 15471 25004 15527 25036
rect 15471 25002 15475 25004
rect 15288 24970 15375 25002
rect 15409 24970 15475 25002
rect 15509 25002 15527 25004
rect 15561 25004 15617 25036
rect 15561 25002 15575 25004
rect 15509 24970 15575 25002
rect 15609 25002 15617 25004
rect 15651 25004 15707 25036
rect 15741 25004 15797 25036
rect 15831 25004 15887 25036
rect 15651 25002 15675 25004
rect 15741 25002 15775 25004
rect 15831 25002 15875 25004
rect 15921 25002 15982 25036
rect 15609 24970 15675 25002
rect 15709 24970 15775 25002
rect 15809 24970 15875 25002
rect 15909 24970 15982 25002
rect 15288 24946 15982 24970
rect 15288 24912 15347 24946
rect 15381 24912 15437 24946
rect 15471 24912 15527 24946
rect 15561 24912 15617 24946
rect 15651 24912 15707 24946
rect 15741 24912 15797 24946
rect 15831 24912 15887 24946
rect 15921 24912 15982 24946
rect 15288 24904 15982 24912
rect 15288 24870 15375 24904
rect 15409 24870 15475 24904
rect 15509 24870 15575 24904
rect 15609 24870 15675 24904
rect 15709 24870 15775 24904
rect 15809 24870 15875 24904
rect 15909 24870 15982 24904
rect 15288 24856 15982 24870
rect 15288 24822 15347 24856
rect 15381 24822 15437 24856
rect 15471 24822 15527 24856
rect 15561 24822 15617 24856
rect 15651 24822 15707 24856
rect 15741 24822 15797 24856
rect 15831 24822 15887 24856
rect 15921 24822 15982 24856
rect 15288 24804 15982 24822
rect 15288 24770 15375 24804
rect 15409 24770 15475 24804
rect 15509 24770 15575 24804
rect 15609 24770 15675 24804
rect 15709 24770 15775 24804
rect 15809 24770 15875 24804
rect 15909 24770 15982 24804
rect 15288 24766 15982 24770
rect 15288 24732 15347 24766
rect 15381 24732 15437 24766
rect 15471 24732 15527 24766
rect 15561 24732 15617 24766
rect 15651 24732 15707 24766
rect 15741 24732 15797 24766
rect 15831 24732 15887 24766
rect 15921 24732 15982 24766
rect 15288 24704 15982 24732
rect 15288 24676 15375 24704
rect 15409 24676 15475 24704
rect 15288 24642 15347 24676
rect 15409 24670 15437 24676
rect 15381 24642 15437 24670
rect 15471 24670 15475 24676
rect 15509 24676 15575 24704
rect 15509 24670 15527 24676
rect 15471 24642 15527 24670
rect 15561 24670 15575 24676
rect 15609 24676 15675 24704
rect 15709 24676 15775 24704
rect 15809 24676 15875 24704
rect 15909 24676 15982 24704
rect 15609 24670 15617 24676
rect 15561 24642 15617 24670
rect 15651 24670 15675 24676
rect 15741 24670 15775 24676
rect 15831 24670 15875 24676
rect 15651 24642 15707 24670
rect 15741 24642 15797 24670
rect 15831 24642 15887 24670
rect 15921 24642 15982 24676
rect 15288 24583 15982 24642
rect 16044 25245 16063 25279
rect 16044 25189 16092 25245
rect 16508 25264 16517 25298
rect 16551 25264 16570 25298
rect 17388 25279 17424 25339
rect 16508 25208 16570 25264
rect 16044 25155 16063 25189
rect 16044 25105 16092 25155
rect 16508 25174 16517 25208
rect 16551 25174 16570 25208
rect 16508 25118 16570 25174
rect 16508 25105 16517 25118
rect 16044 25099 16517 25105
rect 16044 25065 16063 25099
rect 16097 25098 16517 25099
rect 16097 25065 16211 25098
rect 16044 25064 16211 25065
rect 16245 25064 16368 25098
rect 16402 25084 16517 25098
rect 16551 25084 16570 25118
rect 16402 25064 16570 25084
rect 16044 25028 16570 25064
rect 16044 25009 16517 25028
rect 16044 24975 16063 25009
rect 16097 25008 16517 25009
rect 16097 24975 16211 25008
rect 16044 24974 16211 24975
rect 16245 24974 16368 25008
rect 16402 24994 16517 25008
rect 16551 24994 16570 25028
rect 16402 24974 16570 24994
rect 16044 24938 16570 24974
rect 16044 24919 16517 24938
rect 16044 24885 16063 24919
rect 16097 24918 16517 24919
rect 16097 24885 16211 24918
rect 16044 24884 16211 24885
rect 16245 24884 16368 24918
rect 16402 24904 16517 24918
rect 16551 24904 16570 24938
rect 16402 24884 16570 24904
rect 16044 24848 16570 24884
rect 16044 24829 16517 24848
rect 16044 24795 16063 24829
rect 16097 24828 16517 24829
rect 16097 24795 16211 24828
rect 16044 24794 16211 24795
rect 16245 24794 16368 24828
rect 16402 24814 16517 24828
rect 16551 24814 16570 24848
rect 16402 24794 16570 24814
rect 16044 24758 16570 24794
rect 16044 24739 16517 24758
rect 16044 24705 16063 24739
rect 16097 24738 16517 24739
rect 16097 24712 16211 24738
rect 16245 24712 16368 24738
rect 16402 24724 16517 24738
rect 16551 24724 16570 24758
rect 16402 24712 16570 24724
rect 16044 24649 16088 24705
rect 16530 24668 16570 24712
rect 16044 24615 16063 24649
rect 14700 24525 14719 24559
rect 14700 24521 14743 24525
rect 15207 24544 15226 24578
rect 13844 24502 14743 24521
rect 13844 24496 13887 24502
rect 13921 24496 13977 24502
rect 14011 24496 14067 24502
rect 14101 24496 14157 24502
rect 14191 24496 14247 24502
rect 14281 24496 14337 24502
rect 14371 24496 14427 24502
rect 14461 24496 14517 24502
rect 14551 24496 14607 24502
rect 14641 24496 14743 24502
rect 15185 24521 15226 24544
rect 16044 24559 16088 24615
rect 16551 24634 16570 24668
rect 16530 24578 16570 24634
rect 16632 25216 17326 25277
rect 16632 25182 16691 25216
rect 16725 25204 16781 25216
rect 16753 25182 16781 25204
rect 16815 25204 16871 25216
rect 16815 25182 16819 25204
rect 16632 25170 16719 25182
rect 16753 25170 16819 25182
rect 16853 25182 16871 25204
rect 16905 25204 16961 25216
rect 16905 25182 16919 25204
rect 16853 25170 16919 25182
rect 16953 25182 16961 25204
rect 16995 25204 17051 25216
rect 17085 25204 17141 25216
rect 17175 25204 17231 25216
rect 16995 25182 17019 25204
rect 17085 25182 17119 25204
rect 17175 25182 17219 25204
rect 17265 25182 17326 25216
rect 16953 25170 17019 25182
rect 17053 25170 17119 25182
rect 17153 25170 17219 25182
rect 17253 25170 17326 25182
rect 16632 25126 17326 25170
rect 16632 25092 16691 25126
rect 16725 25104 16781 25126
rect 16753 25092 16781 25104
rect 16815 25104 16871 25126
rect 16815 25092 16819 25104
rect 16632 25070 16719 25092
rect 16753 25070 16819 25092
rect 16853 25092 16871 25104
rect 16905 25104 16961 25126
rect 16905 25092 16919 25104
rect 16853 25070 16919 25092
rect 16953 25092 16961 25104
rect 16995 25104 17051 25126
rect 17085 25104 17141 25126
rect 17175 25104 17231 25126
rect 16995 25092 17019 25104
rect 17085 25092 17119 25104
rect 17175 25092 17219 25104
rect 17265 25092 17326 25126
rect 16953 25070 17019 25092
rect 17053 25070 17119 25092
rect 17153 25070 17219 25092
rect 17253 25070 17326 25092
rect 16632 25036 17326 25070
rect 16632 25002 16691 25036
rect 16725 25004 16781 25036
rect 16753 25002 16781 25004
rect 16815 25004 16871 25036
rect 16815 25002 16819 25004
rect 16632 24970 16719 25002
rect 16753 24970 16819 25002
rect 16853 25002 16871 25004
rect 16905 25004 16961 25036
rect 16905 25002 16919 25004
rect 16853 24970 16919 25002
rect 16953 25002 16961 25004
rect 16995 25004 17051 25036
rect 17085 25004 17141 25036
rect 17175 25004 17231 25036
rect 16995 25002 17019 25004
rect 17085 25002 17119 25004
rect 17175 25002 17219 25004
rect 17265 25002 17326 25036
rect 16953 24970 17019 25002
rect 17053 24970 17119 25002
rect 17153 24970 17219 25002
rect 17253 24970 17326 25002
rect 16632 24946 17326 24970
rect 16632 24912 16691 24946
rect 16725 24912 16781 24946
rect 16815 24912 16871 24946
rect 16905 24912 16961 24946
rect 16995 24912 17051 24946
rect 17085 24912 17141 24946
rect 17175 24912 17231 24946
rect 17265 24912 17326 24946
rect 16632 24904 17326 24912
rect 16632 24870 16719 24904
rect 16753 24870 16819 24904
rect 16853 24870 16919 24904
rect 16953 24870 17019 24904
rect 17053 24870 17119 24904
rect 17153 24870 17219 24904
rect 17253 24870 17326 24904
rect 16632 24856 17326 24870
rect 16632 24822 16691 24856
rect 16725 24822 16781 24856
rect 16815 24822 16871 24856
rect 16905 24822 16961 24856
rect 16995 24822 17051 24856
rect 17085 24822 17141 24856
rect 17175 24822 17231 24856
rect 17265 24822 17326 24856
rect 16632 24804 17326 24822
rect 16632 24770 16719 24804
rect 16753 24770 16819 24804
rect 16853 24770 16919 24804
rect 16953 24770 17019 24804
rect 17053 24770 17119 24804
rect 17153 24770 17219 24804
rect 17253 24770 17326 24804
rect 16632 24766 17326 24770
rect 16632 24732 16691 24766
rect 16725 24732 16781 24766
rect 16815 24732 16871 24766
rect 16905 24732 16961 24766
rect 16995 24732 17051 24766
rect 17085 24732 17141 24766
rect 17175 24732 17231 24766
rect 17265 24732 17326 24766
rect 16632 24704 17326 24732
rect 16632 24676 16719 24704
rect 16753 24676 16819 24704
rect 16632 24642 16691 24676
rect 16753 24670 16781 24676
rect 16725 24642 16781 24670
rect 16815 24670 16819 24676
rect 16853 24676 16919 24704
rect 16853 24670 16871 24676
rect 16815 24642 16871 24670
rect 16905 24670 16919 24676
rect 16953 24676 17019 24704
rect 17053 24676 17119 24704
rect 17153 24676 17219 24704
rect 17253 24676 17326 24704
rect 16953 24670 16961 24676
rect 16905 24642 16961 24670
rect 16995 24670 17019 24676
rect 17085 24670 17119 24676
rect 17175 24670 17219 24676
rect 16995 24642 17051 24670
rect 17085 24642 17141 24670
rect 17175 24642 17231 24670
rect 17265 24642 17326 24676
rect 16632 24583 17326 24642
rect 17388 25245 17407 25279
rect 17388 25189 17424 25245
rect 17388 25155 17407 25189
rect 17388 25099 17424 25155
rect 17388 25065 17407 25099
rect 17388 25009 17424 25065
rect 17388 24975 17407 25009
rect 17388 24919 17424 24975
rect 17388 24885 17407 24919
rect 17388 24829 17424 24885
rect 17388 24795 17407 24829
rect 17388 24739 17424 24795
rect 17388 24705 17407 24739
rect 17388 24649 17424 24705
rect 17388 24615 17407 24649
rect 16044 24525 16063 24559
rect 16044 24521 16088 24525
rect 16551 24544 16570 24578
rect 15185 24502 16088 24521
rect 15185 24496 15231 24502
rect 15265 24496 15321 24502
rect 15355 24496 15411 24502
rect 15445 24496 15501 24502
rect 15535 24496 15591 24502
rect 15625 24496 15681 24502
rect 15715 24496 15771 24502
rect 15805 24496 15861 24502
rect 15895 24496 15951 24502
rect 15985 24496 16088 24502
rect 16530 24521 16570 24544
rect 17388 24559 17424 24615
rect 17388 24525 17407 24559
rect 17388 24521 17424 24525
rect 16530 24502 17424 24521
rect 16530 24496 16575 24502
rect 16609 24496 16665 24502
rect 16699 24496 16755 24502
rect 16789 24496 16845 24502
rect 16879 24496 16935 24502
rect 16969 24496 17025 24502
rect 17059 24496 17115 24502
rect 17149 24496 17205 24502
rect 17239 24496 17295 24502
rect 17329 24496 17424 24502
rect 17590 24513 17623 25574
rect 17590 24496 17626 24513
rect 17592 24387 17626 24496
rect 11232 24204 13517 24211
rect 11232 24198 15561 24204
rect 5981 24168 6428 24198
rect 6462 24168 6914 24198
rect 6148 24068 6164 24102
rect 6240 24068 6256 24102
rect 6080 24040 6114 24056
rect 6080 20056 6114 20072
rect 6290 24040 6324 24056
rect 6290 20056 6324 20072
rect 6148 20010 6164 20044
rect 6240 20010 6256 20044
rect 6948 24168 7400 24198
rect 6634 24068 6650 24102
rect 6726 24068 6742 24102
rect 6566 24040 6600 24056
rect 6566 20056 6600 20072
rect 6776 24040 6810 24056
rect 6776 20056 6810 20072
rect 6634 20010 6650 20044
rect 6726 20010 6742 20044
rect 7434 24168 7886 24198
rect 7120 24068 7136 24102
rect 7212 24068 7228 24102
rect 7052 24040 7086 24056
rect 7052 20056 7086 20072
rect 7262 24040 7296 24056
rect 7262 20056 7296 20072
rect 7120 20010 7136 20044
rect 7212 20010 7228 20044
rect 7920 24168 8372 24198
rect 7606 24068 7622 24102
rect 7698 24068 7714 24102
rect 7538 24040 7572 24056
rect 7538 20056 7572 20072
rect 7748 24040 7782 24056
rect 7748 20056 7782 20072
rect 7606 20010 7622 20044
rect 7698 20010 7714 20044
rect 8406 24168 8858 24198
rect 8092 24068 8108 24102
rect 8184 24068 8200 24102
rect 8024 24040 8058 24056
rect 8024 20056 8058 20072
rect 8234 24040 8268 24056
rect 8234 20056 8268 20072
rect 8092 20010 8108 20044
rect 8184 20010 8200 20044
rect 8892 24168 9344 24198
rect 8578 24068 8594 24102
rect 8670 24068 8686 24102
rect 8510 24040 8544 24056
rect 8510 20056 8544 20072
rect 8720 24040 8754 24056
rect 8720 20056 8754 20072
rect 8578 20010 8594 20044
rect 8670 20010 8686 20044
rect 9378 24168 9830 24198
rect 9064 24068 9080 24102
rect 9156 24068 9172 24102
rect 8996 24040 9030 24056
rect 8996 20056 9030 20072
rect 9206 24040 9240 24056
rect 9206 20056 9240 20072
rect 9064 20010 9080 20044
rect 9156 20010 9172 20044
rect 9864 24168 10316 24198
rect 9550 24068 9566 24102
rect 9642 24068 9658 24102
rect 9482 24040 9516 24056
rect 9482 20056 9516 20072
rect 9692 24040 9726 24056
rect 9692 20056 9726 20072
rect 9550 20010 9566 20044
rect 9642 20010 9658 20044
rect 10350 24168 10771 24198
rect 10036 24068 10052 24102
rect 10128 24068 10144 24102
rect 9968 24040 10002 24056
rect 9968 20056 10002 20072
rect 10178 24040 10212 24056
rect 10178 20056 10212 20072
rect 10036 20010 10052 20044
rect 10128 20010 10144 20044
rect 10522 24068 10538 24102
rect 10614 24068 10630 24102
rect 10454 24040 10488 24056
rect 10454 20056 10488 20072
rect 10664 24040 10698 24056
rect 10664 20056 10698 20072
rect 10522 20010 10538 20044
rect 10614 20010 10630 20044
rect 10763 19954 10771 24168
rect 10855 23843 15561 24198
rect 17598 24068 17626 24387
rect 17598 24049 20155 24068
rect 10855 23789 15564 23843
rect 10855 23776 19965 23789
rect 10855 23733 15716 23776
rect 10855 23510 15663 23733
rect 15595 23364 15663 23510
rect 10918 23363 11074 23364
rect 10855 22337 11074 23363
rect 11220 23333 11252 23364
rect 11241 22505 11252 23333
rect 15526 23333 15663 23364
rect 11387 23257 11403 23291
rect 15371 23257 15387 23291
rect 11341 23207 11375 23223
rect 11341 22615 11375 22631
rect 15399 23207 15433 23223
rect 15399 22615 15433 22631
rect 11387 22547 11403 22581
rect 15371 22547 15387 22581
rect 11220 22457 11252 22505
rect 15526 22505 15533 23333
rect 15567 22505 15663 23333
rect 15697 22505 15716 23733
rect 15843 23657 15859 23691
rect 19827 23657 19843 23691
rect 15797 23607 15831 23623
rect 15797 22615 15831 22631
rect 19855 23607 19889 23623
rect 19855 22615 19889 22631
rect 15843 22547 15859 22581
rect 19827 22547 19843 22581
rect 15526 22457 15716 22505
rect 11220 22443 19965 22457
rect 11220 22409 11303 22443
rect 15471 22409 15759 22443
rect 19927 22409 19965 22443
rect 11220 22387 19965 22409
rect 11220 22356 16147 22387
rect 10855 22172 11080 22337
rect 15126 22172 16147 22356
rect 10855 20784 11200 22172
rect 11261 22157 16147 22172
rect 11261 22123 11310 22157
rect 15478 22123 15759 22157
rect 19927 22123 19965 22146
rect 11261 22096 19965 22123
rect 15513 22061 15710 22096
rect 11394 21985 11410 22019
rect 15378 21985 15394 22019
rect 11348 21935 11382 21951
rect 11348 20943 11382 20959
rect 15406 21935 15440 21951
rect 15513 21768 15540 22061
rect 15574 21768 15663 22061
rect 15513 21161 15530 21768
rect 15513 21081 15532 21161
rect 15406 20943 15440 20959
rect 11394 20875 11410 20909
rect 15378 20875 15394 20909
rect 15697 21233 15710 22061
rect 15843 21985 15859 22019
rect 19827 21985 19843 22019
rect 15797 21935 15831 21951
rect 15797 21343 15831 21359
rect 19855 21935 19889 21951
rect 19855 21343 19889 21359
rect 15843 21275 15859 21309
rect 19827 21275 19843 21309
rect 15686 21189 15710 21233
rect 20149 21081 20155 24049
rect 10855 19739 10894 20696
rect 10825 19731 10894 19739
rect 11214 19366 20108 19367
rect 6252 19236 6320 19246
rect 10488 19236 10574 19246
rect 6252 19191 10574 19236
rect 6252 19174 6269 19191
rect 6258 18092 6269 19174
rect 10517 19174 10574 19191
rect 11339 19236 11408 19246
rect 15576 19236 15734 19246
rect 19902 19236 19971 19246
rect 11339 19196 19971 19236
rect 11339 19174 11364 19196
rect 6404 19098 6420 19132
rect 10388 19098 10404 19132
rect 6358 19039 6392 19055
rect 6358 18747 6392 18763
rect 10416 19039 10450 19055
rect 10416 18747 10450 18763
rect 6404 18670 6420 18704
rect 10388 18670 10404 18704
rect 6404 18562 6420 18596
rect 10388 18562 10404 18596
rect 6358 18503 6392 18519
rect 6358 18211 6392 18227
rect 10416 18503 10450 18519
rect 10416 18211 10450 18227
rect 6404 18134 6420 18168
rect 10388 18134 10404 18168
rect 6252 18041 6269 18092
rect 10517 18092 10550 19174
rect 10517 18041 10574 18092
rect 6252 18030 10574 18041
rect 6252 17996 6320 18030
rect 10488 17996 10574 18030
rect 6252 17870 10574 17996
rect 6252 17836 6320 17870
rect 10488 17836 10574 17870
rect 6252 17804 10574 17836
rect 6252 17774 6269 17804
rect 6258 16928 6269 17774
rect 10517 17774 10574 17804
rect 6404 17698 6420 17732
rect 10388 17698 10404 17732
rect 6358 17639 6392 17655
rect 6358 17047 6392 17063
rect 10416 17639 10450 17655
rect 10416 17047 10450 17063
rect 6404 16970 6420 17004
rect 10388 16970 10404 17004
rect 6252 16887 6269 16928
rect 10517 16928 10550 17774
rect 11346 16928 11364 19174
rect 15638 19174 15672 19196
rect 11492 19098 11508 19132
rect 15476 19098 15492 19132
rect 11446 19039 11480 19055
rect 11446 17047 11480 17063
rect 15504 19039 15538 19055
rect 15504 17047 15538 17063
rect 11492 16970 11508 17004
rect 15476 16970 15492 17004
rect 6252 16880 8549 16887
rect 6252 16879 10387 16880
rect 10517 16879 10574 16928
rect 6252 16875 10574 16879
rect 11339 16866 11364 16928
rect 19952 19174 19971 19196
rect 20095 19196 20108 19366
rect 15818 19098 15834 19132
rect 19802 19098 19818 19132
rect 15772 19039 15806 19055
rect 15772 17047 15806 17063
rect 19830 19039 19864 19055
rect 19830 17047 19864 17063
rect 15818 16970 15834 17004
rect 19802 16970 19818 17004
rect 15638 16866 15672 16928
rect 19952 16928 19964 19174
rect 20095 18985 20102 19196
rect 20095 18983 20576 18985
rect 20718 18848 21688 18859
rect 19952 16866 19989 16928
rect 11339 16832 11408 16866
rect 15576 16832 15734 16866
rect 19902 16832 19989 16866
rect 11339 16770 11364 16832
rect 6153 16737 8056 16741
rect 8051 14141 8056 15022
rect 8243 15032 8330 15041
rect 10488 15032 10574 15041
rect 8243 15008 10574 15032
rect 8243 14970 8269 15008
rect 8268 14524 8269 14970
rect 10537 14970 10574 15008
rect 8414 14894 8430 14928
rect 10388 14894 10404 14928
rect 8368 14835 8402 14851
rect 8368 14643 8402 14659
rect 10416 14835 10450 14851
rect 10416 14643 10450 14659
rect 8414 14566 8430 14600
rect 10388 14566 10404 14600
rect 8243 14482 8269 14524
rect 10537 14524 10550 14970
rect 11346 14524 11364 16770
rect 15638 16770 15672 16832
rect 11492 16694 11508 16728
rect 15476 16694 15492 16728
rect 11446 16635 11480 16651
rect 11446 14643 11480 14659
rect 15504 16635 15538 16651
rect 15504 14643 15538 14659
rect 11492 14566 11508 14600
rect 15476 14566 15492 14600
rect 10537 14482 10574 14524
rect 8243 14464 10574 14482
rect 11339 14482 11364 14524
rect 19952 16770 19989 16832
rect 15818 16694 15834 16728
rect 19802 16694 19818 16728
rect 15772 16635 15806 16651
rect 15772 14643 15806 14659
rect 19830 16635 19864 16651
rect 19830 14643 19864 14659
rect 15818 14566 15834 14600
rect 19802 14566 19818 14600
rect 19952 14585 19964 16770
rect 15638 14482 15672 14524
rect 19951 14524 19964 14585
rect 20718 14585 20737 18848
rect 21184 18806 21218 18848
rect 20895 18734 20911 18768
rect 20987 18734 21003 18768
rect 20818 18706 20852 18722
rect 20818 14722 20852 14738
rect 21046 18706 21080 18722
rect 21046 14722 21080 14738
rect 20895 14676 20911 14710
rect 20987 14676 21003 14710
rect 21399 18734 21415 18768
rect 21491 18734 21507 18768
rect 21322 18706 21356 18722
rect 21322 14722 21356 14738
rect 21550 18706 21584 18722
rect 21550 14722 21584 14738
rect 21399 14676 21415 14710
rect 21491 14676 21507 14710
rect 21184 14585 21218 14638
rect 21666 14585 21688 18848
rect 20718 14576 21688 14585
rect 20718 14542 20776 14576
rect 21122 14542 21280 14576
rect 21626 14542 21688 14576
rect 19951 14482 19989 14524
rect 11339 14464 19989 14482
rect 20718 14464 21688 14542
rect 7787 12572 7800 12809
rect 10778 12663 10791 12817
rect 7787 11985 7796 12572
rect 7999 12508 8035 12519
rect 10213 12508 10284 12519
rect 7999 12502 10284 12508
rect 5824 11969 7796 11985
rect 7999 11985 8026 12502
rect 10251 12446 10284 12502
rect 8119 12370 8135 12404
rect 10113 12370 10129 12404
rect 8073 12311 8107 12327
rect 8073 12119 8107 12135
rect 10141 12311 10175 12327
rect 10141 12119 10175 12135
rect 8119 12042 8135 12076
rect 10113 12042 10129 12076
rect 10251 12000 10275 12446
rect 10251 11985 10284 12000
rect 7999 11969 10284 11985
rect 5824 10801 5840 11969
rect 5983 11745 6035 11757
rect 10203 11745 10284 11757
rect 5983 11723 10284 11745
rect 5983 11004 5996 11723
rect 10251 11683 10284 11723
rect 6119 11607 6135 11641
rect 10103 11607 10119 11641
rect 6073 11548 6107 11564
rect 6073 11156 6107 11172
rect 10131 11548 10165 11564
rect 10131 11156 10165 11172
rect 6119 11079 6135 11113
rect 10103 11079 10119 11113
rect 10251 11037 10265 11683
rect 10251 11004 10284 11037
rect 5983 10982 10284 11004
rect 10779 10806 10791 12663
rect 5824 8767 5844 10801
rect 6065 10793 7787 10801
rect 6065 10759 6147 10793
rect 6795 10759 7083 10793
rect 7731 10759 7787 10793
rect 6065 10757 7787 10759
rect 6065 10697 6109 10757
rect 6085 9951 6109 10697
rect 6843 10697 7045 10757
rect 6231 10621 6247 10655
rect 6695 10621 6711 10655
rect 6185 10562 6219 10578
rect 6185 10070 6219 10086
rect 6723 10562 6757 10578
rect 6723 10070 6757 10086
rect 6231 9993 6247 10027
rect 6695 9993 6711 10027
rect 6065 9889 6109 9951
rect 6843 9951 6857 10697
rect 6891 9951 6987 10697
rect 7021 9951 7045 10697
rect 7167 10621 7183 10655
rect 7631 10621 7647 10655
rect 7121 10562 7155 10578
rect 7121 10070 7155 10086
rect 7659 10562 7693 10578
rect 7659 10070 7693 10086
rect 7167 9993 7183 10027
rect 7631 9993 7647 10027
rect 6843 9889 7045 9951
rect 7764 9889 7787 10757
rect 6065 9855 6147 9889
rect 6795 9855 7083 9889
rect 7731 9855 7787 9889
rect 6065 9751 6109 9855
rect 6843 9751 7045 9855
rect 7764 9751 7787 9855
rect 6065 9717 6147 9751
rect 6795 9717 7083 9751
rect 7731 9717 7787 9751
rect 6065 9655 6109 9717
rect 6085 8909 6109 9655
rect 6843 9655 7045 9717
rect 6231 9579 6247 9613
rect 6695 9579 6711 9613
rect 6185 9520 6219 9536
rect 6185 9028 6219 9044
rect 6723 9520 6757 9536
rect 6723 9028 6757 9044
rect 6231 8951 6247 8985
rect 6695 8951 6711 8985
rect 6065 8884 6109 8909
rect 6843 8909 6857 9655
rect 6891 8909 6987 9655
rect 7021 8909 7045 9655
rect 7167 9579 7183 9613
rect 7631 9579 7647 9613
rect 7121 9520 7155 9536
rect 7121 9028 7155 9044
rect 7659 9520 7693 9536
rect 7659 9028 7693 9044
rect 7167 8951 7183 8985
rect 7631 8951 7647 8985
rect 6843 8884 7045 8909
rect 7764 8884 7787 9717
rect 6065 8871 7787 8884
rect 7942 8871 8812 10801
rect 8950 10777 9013 10801
rect 9661 10777 9945 10801
rect 10593 10777 10655 10806
rect 8950 10757 10655 10777
rect 8950 10715 8978 10757
rect 8951 9969 8978 10715
rect 9721 10715 9905 10757
rect 9097 10639 9113 10673
rect 9561 10639 9577 10673
rect 9051 10580 9085 10596
rect 9051 10088 9085 10104
rect 9589 10580 9623 10596
rect 9589 10088 9623 10104
rect 9097 10011 9113 10045
rect 9561 10011 9577 10045
rect 8950 9936 8978 9969
rect 9721 9969 9723 10715
rect 9757 9969 9849 10715
rect 9883 9969 9905 10715
rect 10029 10639 10045 10673
rect 10493 10639 10509 10673
rect 9983 10580 10017 10596
rect 9983 10088 10017 10104
rect 10521 10580 10555 10596
rect 10521 10088 10555 10104
rect 10029 10011 10045 10045
rect 10493 10011 10509 10045
rect 9721 9936 9905 9969
rect 10633 9936 10655 10757
rect 8950 9907 10655 9936
rect 8950 9873 9013 9907
rect 9661 9873 9945 9907
rect 10593 9873 10655 9907
rect 8950 9726 10655 9873
rect 8950 9692 9013 9726
rect 9661 9692 9945 9726
rect 10593 9692 10655 9726
rect 8950 9684 10655 9692
rect 8950 9630 8978 9684
rect 8951 8884 8978 9630
rect 9721 9630 9905 9684
rect 9097 9554 9113 9588
rect 9561 9554 9577 9588
rect 9051 9495 9085 9511
rect 9051 9003 9085 9019
rect 9589 9495 9623 9511
rect 9589 9003 9623 9019
rect 9097 8926 9113 8960
rect 9561 8926 9577 8960
rect 9721 8884 9723 9630
rect 9757 8884 9849 9630
rect 9883 8884 9905 9630
rect 10029 9554 10045 9588
rect 10493 9554 10509 9588
rect 9983 9495 10017 9511
rect 9983 9003 10017 9019
rect 10521 9495 10555 9511
rect 10521 9003 10555 9019
rect 10029 8926 10045 8960
rect 10493 8926 10509 8960
rect 7960 8767 8812 8871
rect 8950 8877 9015 8884
rect 9721 8877 9905 8884
rect 10633 8877 10655 9684
rect 8950 8863 10655 8877
rect 5824 8749 8812 8767
rect 5824 8742 6109 8749
rect 10776 8742 10791 10806
rect 11839 11117 12918 11128
rect 11839 11114 11880 11117
rect 11839 10511 11848 11114
rect 12899 11079 12918 11117
rect 11967 10991 12773 11006
rect 11836 10404 11848 10511
rect 11967 10511 11994 10991
rect 12079 10912 12095 10946
rect 12163 10912 12179 10946
rect 12237 10912 12253 10946
rect 12321 10912 12337 10946
rect 12395 10912 12411 10946
rect 12479 10912 12495 10946
rect 12553 10912 12569 10946
rect 12637 10912 12653 10946
rect 12033 10853 12067 10869
rect 12033 10661 12067 10677
rect 12191 10853 12225 10869
rect 12191 10661 12225 10677
rect 12349 10853 12383 10869
rect 12349 10661 12383 10677
rect 12507 10853 12541 10869
rect 12507 10661 12541 10677
rect 12665 10853 12699 10869
rect 12665 10661 12699 10677
rect 12079 10584 12095 10618
rect 12163 10584 12179 10618
rect 12237 10584 12253 10618
rect 12321 10584 12337 10618
rect 12395 10584 12411 10618
rect 12479 10584 12495 10618
rect 12553 10584 12569 10618
rect 12637 10584 12653 10618
rect 12763 10511 12773 10991
rect 11967 10507 12773 10511
rect 11967 10473 11973 10507
rect 12757 10473 12773 10507
rect 11967 10418 12773 10473
rect 12901 10418 12918 11079
rect 13691 11042 20445 11076
rect 13691 10789 13753 11042
rect 20417 10853 20445 11042
rect 11967 10404 12918 10418
rect 11836 10352 12918 10404
rect 11228 9901 13466 9915
rect 11228 9898 12280 9901
rect 11228 9173 11241 9898
rect 11310 9860 11723 9898
rect 11310 9826 11379 9860
rect 11647 9826 11723 9860
rect 11310 9764 11329 9826
rect 11317 9336 11329 9764
rect 11709 9764 11723 9826
rect 11848 9860 12280 9898
rect 11848 9826 11935 9860
rect 12203 9826 12280 9860
rect 11848 9764 11873 9826
rect 11463 9688 11479 9722
rect 11547 9688 11563 9722
rect 11417 9638 11451 9654
rect 11417 9446 11451 9462
rect 11575 9638 11609 9654
rect 11575 9446 11609 9462
rect 11463 9378 11479 9412
rect 11547 9378 11563 9412
rect 11310 9301 11329 9336
rect 12265 9764 12280 9826
rect 12405 9900 13466 9901
rect 12405 9893 13384 9900
rect 12405 9860 12844 9893
rect 12405 9826 12491 9860
rect 12759 9826 12844 9860
rect 12405 9764 12429 9826
rect 12019 9688 12035 9722
rect 12103 9688 12119 9722
rect 11973 9638 12007 9654
rect 11973 9446 12007 9462
rect 12131 9638 12165 9654
rect 12131 9446 12165 9462
rect 12019 9378 12035 9412
rect 12103 9378 12119 9412
rect 11709 9301 11723 9336
rect 11310 9287 11723 9301
rect 11848 9301 11873 9336
rect 12820 9764 12844 9826
rect 12969 9860 13384 9893
rect 12969 9826 13047 9860
rect 13315 9826 13384 9860
rect 12969 9764 12985 9826
rect 12575 9688 12591 9722
rect 12659 9688 12675 9722
rect 12529 9638 12563 9654
rect 12529 9446 12563 9462
rect 12687 9638 12721 9654
rect 12687 9446 12721 9462
rect 12575 9378 12591 9412
rect 12659 9378 12675 9412
rect 12265 9301 12280 9336
rect 11848 9287 12280 9301
rect 12405 9301 12429 9336
rect 12820 9336 12821 9764
rect 13375 9764 13384 9826
rect 13131 9688 13147 9722
rect 13215 9688 13231 9722
rect 13085 9638 13119 9654
rect 13085 9446 13119 9462
rect 13243 9638 13277 9654
rect 13243 9446 13277 9462
rect 13131 9378 13147 9412
rect 13215 9378 13231 9412
rect 12820 9301 12844 9336
rect 12405 9287 12844 9301
rect 12969 9301 12985 9336
rect 13375 9336 13377 9764
rect 13375 9301 13384 9336
rect 12969 9287 13384 9301
rect 13448 9287 13466 9900
rect 13446 9173 13466 9287
rect 11228 9141 13466 9173
rect 6828 8651 7060 8655
rect 8924 8651 10822 8655
rect 5282 8650 10822 8651
rect 5282 8640 8523 8650
rect 5282 8630 5318 8640
rect 5282 5730 5295 8630
rect 8589 8626 10822 8650
rect 5375 8543 8523 8560
rect 5375 8045 5390 8543
rect 6828 8513 7060 8543
rect 5511 8437 5527 8471
rect 6695 8437 6711 8471
rect 5465 8387 5499 8403
rect 5465 8195 5499 8211
rect 6723 8387 6757 8403
rect 6723 8195 6757 8211
rect 5511 8127 5527 8161
rect 6695 8127 6711 8161
rect 6828 8085 6857 8513
rect 6891 8085 6987 8513
rect 7021 8085 7060 8513
rect 8495 8513 8523 8543
rect 7167 8437 7183 8471
rect 8351 8437 8367 8471
rect 7121 8387 7155 8403
rect 7121 8195 7155 8211
rect 8379 8387 8413 8403
rect 8379 8195 8413 8211
rect 7167 8127 7183 8161
rect 8351 8127 8367 8161
rect 6828 8045 7060 8085
rect 8495 8085 8513 8513
rect 8495 8045 8523 8085
rect 5375 8023 8523 8045
rect 5375 8009 5427 8023
rect 6795 8009 7083 8023
rect 8451 8009 8523 8023
rect 8589 7995 8824 8564
rect 8961 8539 9704 8564
rect 8961 8058 8967 8539
rect 9654 8513 9704 8539
rect 9897 8539 10665 8564
rect 9897 8514 9955 8539
rect 9097 8437 9113 8471
rect 9521 8437 9537 8471
rect 9051 8387 9085 8403
rect 9051 8195 9085 8211
rect 9549 8387 9583 8403
rect 9549 8195 9583 8211
rect 9097 8127 9113 8161
rect 9521 8127 9537 8161
rect 9654 8085 9683 8513
rect 9923 8086 9955 8514
rect 10637 8514 10665 8539
rect 10069 8438 10085 8472
rect 10493 8438 10509 8472
rect 10023 8388 10057 8404
rect 10023 8196 10057 8212
rect 10521 8388 10555 8404
rect 10521 8196 10555 8212
rect 10069 8128 10085 8162
rect 10493 8128 10509 8162
rect 9654 8058 9704 8085
rect 8961 8023 9704 8058
rect 8961 7995 9013 8023
rect 9621 7995 9704 8023
rect 9897 8058 9955 8086
rect 10637 8086 10655 8514
rect 10637 8058 10665 8086
rect 9897 8024 10665 8058
rect 9897 7995 9985 8024
rect 10593 7995 10665 8024
rect 10790 8058 10822 8626
rect 10790 7995 10826 8058
rect 10802 7933 10826 7995
rect 8589 7891 10826 7933
rect 5375 7859 5427 7869
rect 6795 7859 7083 7869
rect 8451 7859 8523 7869
rect 5375 7836 8523 7859
rect 5375 7334 5390 7836
rect 6828 7797 7060 7836
rect 5511 7721 5527 7755
rect 6695 7721 6711 7755
rect 5465 7671 5499 7687
rect 5465 7479 5499 7495
rect 6723 7671 6757 7687
rect 6723 7479 6757 7495
rect 5511 7411 5527 7445
rect 6695 7411 6711 7445
rect 6828 7369 6857 7797
rect 6891 7369 6987 7797
rect 7021 7369 7060 7797
rect 8495 7797 8523 7836
rect 7167 7721 7183 7755
rect 8351 7721 8367 7755
rect 7121 7671 7155 7687
rect 7121 7479 7155 7495
rect 8379 7671 8413 7687
rect 8379 7479 8413 7495
rect 7167 7411 7183 7445
rect 8351 7411 8367 7445
rect 6828 7334 7060 7369
rect 8495 7369 8513 7797
rect 8495 7334 8523 7369
rect 5375 7307 8523 7334
rect 5375 7295 5427 7307
rect 6795 7295 7083 7307
rect 8451 7295 8523 7307
rect 5375 7143 5427 7155
rect 6795 7143 7083 7155
rect 8451 7143 8523 7155
rect 5375 7125 8523 7143
rect 5375 6610 5390 7125
rect 6828 7081 7060 7125
rect 5511 7005 5527 7039
rect 6695 7005 6711 7039
rect 5465 6955 5499 6971
rect 5465 6763 5499 6779
rect 6723 6955 6757 6971
rect 6723 6763 6757 6779
rect 5511 6695 5527 6729
rect 6695 6695 6711 6729
rect 6828 6653 6857 7081
rect 6891 6653 6987 7081
rect 7021 6653 7060 7081
rect 8495 7081 8523 7125
rect 7167 7005 7183 7039
rect 8351 7005 8367 7039
rect 7121 6955 7155 6971
rect 7121 6763 7155 6779
rect 8379 6955 8413 6971
rect 8379 6763 8413 6779
rect 7167 6695 7183 6729
rect 8351 6695 8367 6729
rect 6828 6610 7060 6653
rect 8495 6653 8513 7081
rect 8495 6610 8523 6653
rect 5375 6591 8523 6610
rect 5375 6564 5427 6591
rect 6795 6564 7083 6591
rect 8451 6564 8523 6591
rect 5375 6401 8523 6424
rect 5375 5911 5390 6401
rect 6828 6365 7060 6401
rect 5511 6289 5527 6323
rect 6695 6289 6711 6323
rect 5465 6239 5499 6255
rect 5465 6047 5499 6063
rect 6723 6239 6757 6255
rect 6723 6047 6757 6063
rect 5511 5979 5527 6013
rect 6695 5979 6711 6013
rect 6828 5937 6857 6365
rect 6891 5937 6987 6365
rect 7021 5937 7060 6365
rect 8495 6365 8523 6401
rect 7167 6289 7183 6323
rect 8351 6289 8367 6323
rect 7121 6239 7155 6255
rect 7121 6047 7155 6063
rect 8379 6239 8413 6255
rect 8379 6047 8413 6063
rect 7167 5979 7183 6013
rect 8351 5979 8367 6013
rect 6828 5911 7060 5937
rect 8495 5937 8513 6365
rect 8495 5911 8523 5937
rect 5375 5875 8523 5911
rect 5375 5867 5427 5875
rect 6795 5867 7083 5875
rect 8451 5867 8523 5875
rect 5282 5727 5335 5730
rect 5282 5720 8523 5727
rect 8589 5720 8632 7891
rect 10637 7886 10822 7891
rect 5282 5709 8632 5720
rect 8495 5705 8632 5709
rect 13692 2259 13753 10789
rect 13873 10827 20445 10853
rect 13873 10793 14063 10827
rect 14201 10793 14359 10827
rect 14497 10793 14655 10827
rect 14793 10793 14951 10827
rect 15089 10793 15247 10827
rect 15385 10793 15543 10827
rect 15681 10793 15839 10827
rect 15977 10793 16135 10827
rect 16273 10793 20445 10827
rect 13873 10789 20445 10793
rect 13873 10731 14009 10789
rect 13873 6731 13967 10731
rect 14001 6731 14009 10731
rect 14263 10731 14297 10789
rect 13873 6669 14009 6731
rect 14559 10731 14593 10789
rect 14263 6669 14297 6731
rect 14855 10731 14889 10789
rect 14559 6669 14593 6731
rect 15151 10731 15185 10789
rect 14855 6669 14889 6731
rect 15447 10731 15481 10789
rect 15151 6669 15185 6731
rect 15743 10731 15777 10789
rect 15447 6669 15481 6731
rect 16039 10731 16073 10789
rect 15743 6669 15777 6731
rect 16330 10731 20445 10789
rect 16330 9873 16335 10731
rect 16039 6669 16073 6731
rect 16318 6731 16335 9873
rect 16369 10288 20445 10731
rect 16369 10100 16585 10288
rect 20388 10277 20445 10288
rect 16369 9898 20274 10100
rect 16369 9864 16571 9898
rect 20157 9864 20274 9898
rect 16369 9830 20274 9864
rect 16369 9802 16544 9830
rect 16369 7574 16475 9802
rect 16509 7574 16544 9802
rect 20197 9802 20274 9830
rect 16655 9726 16671 9760
rect 16739 9726 16755 9760
rect 16813 9726 16829 9760
rect 16897 9726 16913 9760
rect 16971 9726 16987 9760
rect 17055 9726 17071 9760
rect 17129 9726 17145 9760
rect 17213 9726 17229 9760
rect 17287 9726 17303 9760
rect 17371 9726 17387 9760
rect 17445 9726 17461 9760
rect 17529 9726 17545 9760
rect 17603 9726 17619 9760
rect 17687 9726 17703 9760
rect 17761 9726 17777 9760
rect 17845 9726 17861 9760
rect 17919 9726 17935 9760
rect 18003 9726 18019 9760
rect 18077 9726 18093 9760
rect 18161 9726 18177 9760
rect 18235 9726 18251 9760
rect 18319 9726 18335 9760
rect 18393 9726 18409 9760
rect 18477 9726 18493 9760
rect 18551 9726 18567 9760
rect 18635 9726 18651 9760
rect 18709 9726 18725 9760
rect 18793 9726 18809 9760
rect 18867 9726 18883 9760
rect 18951 9726 18967 9760
rect 19025 9726 19041 9760
rect 19109 9726 19125 9760
rect 19183 9726 19199 9760
rect 19267 9726 19283 9760
rect 19341 9726 19357 9760
rect 19425 9726 19441 9760
rect 19499 9726 19515 9760
rect 19583 9726 19599 9760
rect 19657 9726 19673 9760
rect 19741 9726 19757 9760
rect 19815 9726 19831 9760
rect 19899 9726 19915 9760
rect 19973 9726 19989 9760
rect 20057 9726 20073 9760
rect 16609 9676 16643 9692
rect 16609 7684 16643 7700
rect 16767 9676 16801 9692
rect 16767 7684 16801 7700
rect 16925 9676 16959 9692
rect 16925 7684 16959 7700
rect 17083 9676 17117 9692
rect 17083 7684 17117 7700
rect 17241 9676 17275 9692
rect 17241 7684 17275 7700
rect 17399 9676 17433 9692
rect 17399 7684 17433 7700
rect 17557 9676 17591 9692
rect 17557 7684 17591 7700
rect 17715 9676 17749 9692
rect 17715 7684 17749 7700
rect 17873 9676 17907 9692
rect 17873 7684 17907 7700
rect 18031 9676 18065 9692
rect 18031 7684 18065 7700
rect 18189 9676 18223 9692
rect 18189 7684 18223 7700
rect 18347 9676 18381 9692
rect 18347 7684 18381 7700
rect 18505 9676 18539 9692
rect 18505 7684 18539 7700
rect 18663 9676 18697 9692
rect 18663 7684 18697 7700
rect 18821 9676 18855 9692
rect 18821 7684 18855 7700
rect 18979 9676 19013 9692
rect 18979 7684 19013 7700
rect 19137 9676 19171 9692
rect 19137 7684 19171 7700
rect 19295 9676 19329 9692
rect 19295 7684 19329 7700
rect 19453 9676 19487 9692
rect 19453 7684 19487 7700
rect 19611 9676 19645 9692
rect 19611 7684 19645 7700
rect 19769 9676 19803 9692
rect 19769 7684 19803 7700
rect 19927 9676 19961 9692
rect 19927 7684 19961 7700
rect 20085 9676 20119 9692
rect 20085 7684 20119 7700
rect 16655 7616 16671 7650
rect 16739 7616 16755 7650
rect 16813 7616 16829 7650
rect 16897 7616 16913 7650
rect 16971 7616 16987 7650
rect 17055 7616 17071 7650
rect 17129 7616 17145 7650
rect 17213 7616 17229 7650
rect 17287 7616 17303 7650
rect 17371 7616 17387 7650
rect 17445 7616 17461 7650
rect 17529 7616 17545 7650
rect 17603 7616 17619 7650
rect 17687 7616 17703 7650
rect 17761 7616 17777 7650
rect 17845 7616 17861 7650
rect 17919 7616 17935 7650
rect 18003 7616 18019 7650
rect 18077 7616 18093 7650
rect 18161 7616 18177 7650
rect 18235 7616 18251 7650
rect 18319 7616 18335 7650
rect 18393 7616 18409 7650
rect 18477 7616 18493 7650
rect 18551 7616 18567 7650
rect 18635 7616 18651 7650
rect 18709 7616 18725 7650
rect 18793 7616 18809 7650
rect 18867 7616 18883 7650
rect 18951 7616 18967 7650
rect 19025 7616 19041 7650
rect 19109 7616 19125 7650
rect 19183 7616 19199 7650
rect 19267 7616 19283 7650
rect 19341 7616 19357 7650
rect 19425 7616 19441 7650
rect 19499 7616 19515 7650
rect 19583 7616 19599 7650
rect 19657 7616 19673 7650
rect 19741 7616 19757 7650
rect 19815 7616 19831 7650
rect 19899 7616 19915 7650
rect 19973 7616 19989 7650
rect 20057 7616 20073 7650
rect 16369 7533 16544 7574
rect 20197 7574 20219 9802
rect 20253 7574 20274 9802
rect 20197 7533 20274 7574
rect 16369 7512 20274 7533
rect 16369 7478 16571 7512
rect 20157 7478 20274 7512
rect 16369 7473 20274 7478
rect 16369 7290 16471 7473
rect 16369 7277 16567 7290
rect 16995 7277 17153 7290
rect 17581 7277 17739 7290
rect 18167 7277 20160 7290
rect 16369 7264 20160 7277
rect 16369 7215 16544 7264
rect 16369 6731 16471 7215
rect 16318 6669 16471 6731
rect 13873 6635 14063 6669
rect 14201 6635 14359 6669
rect 14497 6635 14655 6669
rect 14793 6635 14951 6669
rect 15089 6635 15247 6669
rect 15385 6635 15543 6669
rect 15681 6635 15839 6669
rect 15977 6635 16135 6669
rect 16273 6635 16471 6669
rect 13873 6573 14009 6635
rect 13873 2573 13967 6573
rect 14001 2573 14009 6573
rect 14263 6573 14297 6635
rect 13873 2540 14009 2573
rect 14559 6573 14593 6635
rect 14263 2540 14297 2573
rect 14855 6573 14889 6635
rect 14559 2540 14593 2573
rect 15151 6573 15185 6635
rect 14855 2540 14889 2573
rect 15447 6573 15481 6635
rect 15151 2540 15185 2573
rect 15743 6573 15777 6635
rect 15447 2540 15481 2573
rect 16039 6573 16073 6635
rect 15743 2540 15777 2573
rect 16318 6573 16471 6635
rect 16039 2540 16073 2573
rect 16318 2573 16335 6573
rect 16369 5047 16471 6573
rect 16505 5047 16544 7215
rect 17057 7215 17091 7264
rect 16677 7143 16693 7177
rect 16869 7143 16885 7177
rect 16609 7115 16643 7131
rect 16609 5131 16643 5147
rect 16919 7115 16953 7131
rect 16919 5131 16953 5147
rect 16677 5085 16693 5119
rect 16869 5085 16885 5119
rect 16369 4985 16544 5047
rect 17643 7215 17677 7264
rect 17263 7143 17279 7177
rect 17455 7143 17471 7177
rect 17195 7115 17229 7131
rect 17195 5131 17229 5147
rect 17505 7115 17539 7131
rect 17505 5131 17539 5147
rect 17263 5085 17279 5119
rect 17455 5085 17471 5119
rect 17057 4985 17091 5047
rect 18229 7215 20160 7264
rect 17849 7143 17865 7177
rect 18041 7143 18057 7177
rect 17781 7115 17815 7131
rect 17781 5131 17815 5147
rect 18091 7115 18125 7131
rect 18091 5131 18125 5147
rect 17849 5085 17865 5119
rect 18041 5085 18057 5119
rect 17643 4985 17677 5047
rect 18263 6561 20160 7215
rect 18263 6378 18519 6561
rect 19526 6378 20160 6561
rect 18263 6369 20160 6378
rect 18263 6335 18680 6369
rect 18818 6335 18976 6369
rect 19114 6335 19272 6369
rect 19410 6335 19568 6369
rect 19706 6335 20160 6369
rect 18263 6330 20160 6335
rect 18263 6273 18621 6330
rect 18263 5047 18584 6273
rect 18229 4985 18584 5047
rect 16369 4951 16567 4985
rect 16995 4951 17153 4985
rect 17581 4951 17739 4985
rect 18167 4951 18584 4985
rect 16369 4849 16544 4951
rect 18236 4849 18584 4951
rect 16369 4815 16567 4849
rect 16995 4815 17153 4849
rect 17581 4815 17739 4849
rect 18167 4815 18584 4849
rect 16369 4753 16544 4815
rect 16369 2585 16471 4753
rect 16505 2585 16544 4753
rect 17057 4753 17091 4815
rect 16677 4681 16693 4715
rect 16869 4681 16885 4715
rect 16609 4653 16643 4669
rect 16609 2669 16643 2685
rect 16919 4653 16953 4669
rect 16919 2669 16953 2685
rect 16677 2623 16693 2657
rect 16869 2623 16885 2657
rect 16369 2573 16544 2585
rect 16318 2540 16544 2573
rect 17643 4753 17677 4815
rect 17263 4681 17279 4715
rect 17455 4681 17471 4715
rect 17195 4653 17229 4669
rect 17195 2669 17229 2685
rect 17505 4653 17539 4669
rect 17505 2669 17539 2685
rect 17263 2623 17279 2657
rect 17455 2623 17471 2657
rect 17057 2540 17091 2585
rect 18229 4753 18584 4815
rect 17849 4681 17865 4715
rect 18041 4681 18057 4715
rect 17781 4653 17815 4669
rect 17781 2669 17815 2685
rect 18091 4653 18125 4669
rect 18091 2669 18125 2685
rect 17849 2623 17865 2657
rect 18041 2623 18057 2657
rect 17643 2540 17677 2585
rect 18263 2585 18584 4753
rect 18229 2573 18584 2585
rect 18618 2573 18621 6273
rect 18880 6273 18914 6330
rect 18229 2540 18621 2573
rect 19176 6273 19210 6330
rect 18880 2540 18914 2573
rect 19472 6273 19506 6330
rect 19176 2540 19210 2573
rect 19768 6273 20160 6330
rect 19472 2540 19506 2573
rect 19802 2573 20160 6273
rect 19768 2540 20160 2573
rect 13873 2523 20160 2540
rect 13873 2511 16567 2523
rect 13873 2477 14063 2511
rect 14201 2477 14359 2511
rect 14497 2477 14655 2511
rect 14793 2477 14951 2511
rect 15089 2477 15247 2511
rect 15385 2477 15543 2511
rect 15681 2477 15839 2511
rect 15977 2477 16135 2511
rect 16273 2489 16567 2511
rect 16995 2489 17153 2523
rect 17581 2489 17739 2523
rect 18167 2511 20160 2523
rect 18167 2489 18680 2511
rect 16273 2477 18680 2489
rect 18818 2477 18976 2511
rect 19114 2477 19272 2511
rect 19410 2477 19568 2511
rect 19706 2477 20160 2511
rect 13873 2391 20160 2477
rect 13692 2254 20160 2259
rect 20400 2254 20445 10277
rect 13692 2211 20445 2254
rect 21186 8161 24142 8179
rect 21186 8145 21325 8161
rect 21186 3233 21195 8145
rect 24025 8129 24142 8161
rect 21504 7988 23911 8031
rect 21504 7983 21585 7988
rect 21504 6015 21527 7983
rect 21561 6015 21585 7983
rect 21733 7911 21749 7945
rect 23725 7911 23741 7945
rect 21665 7883 21699 7899
rect 21665 6099 21699 6115
rect 23775 7883 23809 7899
rect 23775 6099 23809 6115
rect 21733 6053 21749 6087
rect 23725 6053 23741 6087
rect 21504 5971 21585 6015
rect 23885 5971 23911 7988
rect 21504 5964 23911 5971
rect 23723 5953 23911 5964
rect 23851 5919 23911 5953
rect 23723 5829 23911 5919
rect 23851 5795 23911 5829
rect 21504 5788 23911 5795
rect 21504 5733 21585 5788
rect 21504 3765 21527 5733
rect 21561 3765 21585 5733
rect 21733 5661 21749 5695
rect 23725 5661 23741 5695
rect 21665 5633 21699 5649
rect 21665 3849 21699 3865
rect 23775 5633 23809 5649
rect 23775 3849 23809 3865
rect 23885 4060 23911 5788
rect 24090 4362 24142 8129
rect 24321 8168 26867 8179
rect 24321 7835 24363 8168
rect 25879 8159 26867 8168
rect 26789 8149 26867 8159
rect 24619 8034 25836 8040
rect 24619 7983 24689 8034
rect 24321 5025 24364 7835
rect 24646 7615 24689 7983
rect 25801 7983 25836 8034
rect 24827 7911 24843 7945
rect 25619 7911 25635 7945
rect 24750 7883 24784 7899
rect 24750 7699 24784 7715
rect 25678 7883 25712 7899
rect 25678 7699 25712 7715
rect 24827 7653 24843 7687
rect 25619 7653 25635 7687
rect 24618 7567 24689 7615
rect 25801 7615 25816 7983
rect 25801 7567 25836 7615
rect 24618 7553 25836 7567
rect 24618 7519 24708 7553
rect 25754 7537 25836 7553
rect 24618 7373 24883 7519
rect 24618 7339 24708 7373
rect 26654 7339 26708 7369
rect 24618 7317 26708 7339
rect 24618 7277 24689 7317
rect 24646 5103 24689 7277
rect 24827 7205 24843 7239
rect 26519 7205 26535 7239
rect 24750 7177 24784 7193
rect 24750 6993 24784 7009
rect 26578 7177 26612 7193
rect 26578 6993 26612 7009
rect 24827 6947 24843 6981
rect 26519 6947 26535 6981
rect 24750 6919 24784 6935
rect 24750 6735 24784 6751
rect 26578 6919 26612 6935
rect 26578 6735 26612 6751
rect 24827 6689 24843 6723
rect 26519 6689 26535 6723
rect 24750 6661 24784 6677
rect 24750 6477 24784 6493
rect 26578 6661 26612 6677
rect 26578 6477 26612 6493
rect 24827 6431 24843 6465
rect 26519 6431 26535 6465
rect 24750 6403 24784 6419
rect 24750 6219 24784 6235
rect 26578 6403 26612 6419
rect 26578 6219 26612 6235
rect 24827 6173 24843 6207
rect 26519 6173 26535 6207
rect 24750 6145 24784 6161
rect 24750 5961 24784 5977
rect 26578 6145 26612 6161
rect 26578 5961 26612 5977
rect 24827 5915 24843 5949
rect 26519 5915 26535 5949
rect 24750 5887 24784 5903
rect 24750 5703 24784 5719
rect 26578 5887 26612 5903
rect 26578 5703 26612 5719
rect 24827 5657 24843 5691
rect 26519 5657 26535 5691
rect 24750 5629 24784 5645
rect 24750 5445 24784 5461
rect 26578 5629 26612 5645
rect 26578 5445 26612 5461
rect 24827 5399 24843 5433
rect 26519 5399 26535 5433
rect 24750 5371 24784 5387
rect 24750 5187 24784 5203
rect 26578 5371 26612 5387
rect 26578 5187 26612 5203
rect 24827 5141 24843 5175
rect 26519 5141 26535 5175
rect 24618 5081 24689 5103
rect 26669 5081 26708 7317
rect 24618 5041 26708 5081
rect 24618 5025 24708 5041
rect 26654 5025 26708 5041
rect 24321 4469 24358 5025
rect 26835 4469 26867 8149
rect 24321 4449 26867 4469
rect 24090 4311 26918 4362
rect 21733 3803 21749 3837
rect 23725 3803 23741 3837
rect 21504 3725 21585 3765
rect 23885 3765 23913 4060
rect 23947 4050 24020 4060
rect 23947 3971 26830 4050
rect 23947 3937 24552 3971
rect 26780 3937 26830 3971
rect 23947 3875 24528 3937
rect 23947 3765 24456 3875
rect 23885 3744 24456 3765
rect 23885 3725 23911 3744
rect 21504 3703 23911 3725
rect 21504 3669 21623 3703
rect 23851 3669 23911 3703
rect 21504 3591 23911 3669
rect 24090 3591 24456 3744
rect 21186 1656 21199 3233
rect 24301 3201 24456 3591
rect 24290 3147 24456 3201
rect 21328 3103 21408 3106
rect 24098 3103 24187 3106
rect 21328 3083 24187 3103
rect 21328 3041 21362 3083
rect 21346 1813 21362 3041
rect 24150 3041 24187 3083
rect 21492 2965 21508 2999
rect 21676 2965 21692 2999
rect 21750 2965 21766 2999
rect 21934 2965 21950 2999
rect 22008 2965 22024 2999
rect 22192 2965 22208 2999
rect 22266 2965 22282 2999
rect 22450 2965 22466 2999
rect 22524 2965 22540 2999
rect 22708 2965 22724 2999
rect 22782 2965 22798 2999
rect 22966 2965 22982 2999
rect 23040 2965 23056 2999
rect 23224 2965 23240 2999
rect 23298 2965 23314 2999
rect 23482 2965 23498 2999
rect 23556 2965 23572 2999
rect 23740 2965 23756 2999
rect 23814 2965 23830 2999
rect 23998 2965 24014 2999
rect 21446 2915 21480 2931
rect 21446 1923 21480 1939
rect 21704 2915 21738 2931
rect 21704 1923 21738 1939
rect 21962 2915 21996 2931
rect 21962 1923 21996 1939
rect 22220 2915 22254 2931
rect 22220 1923 22254 1939
rect 22478 2915 22512 2931
rect 22478 1923 22512 1939
rect 22736 2915 22770 2931
rect 22736 1923 22770 1939
rect 22994 2915 23028 2931
rect 22994 1923 23028 1939
rect 23252 2915 23286 2931
rect 23252 1923 23286 1939
rect 23510 2915 23544 2931
rect 23510 1923 23544 1939
rect 23768 2915 23802 2931
rect 23768 1923 23802 1939
rect 24026 2915 24060 2931
rect 24026 1923 24060 1939
rect 21492 1855 21508 1889
rect 21676 1855 21692 1889
rect 21750 1855 21766 1889
rect 21934 1855 21950 1889
rect 22008 1855 22024 1889
rect 22192 1855 22208 1889
rect 22266 1855 22282 1889
rect 22450 1855 22466 1889
rect 22524 1855 22540 1889
rect 22708 1855 22724 1889
rect 22782 1855 22798 1889
rect 22966 1855 22982 1889
rect 23040 1855 23056 1889
rect 23224 1855 23240 1889
rect 23298 1855 23314 1889
rect 23482 1855 23498 1889
rect 23556 1855 23572 1889
rect 23740 1855 23756 1889
rect 23814 1855 23830 1889
rect 23998 1855 24014 1889
rect 21328 1805 21362 1813
rect 24150 1813 24160 3041
rect 24295 1907 24456 3147
rect 24490 1907 24528 3875
rect 24662 3803 24678 3837
rect 26654 3803 26670 3837
rect 24594 3775 24628 3791
rect 24594 1991 24628 2007
rect 26704 3775 26738 3791
rect 26704 1991 26738 2007
rect 24662 1945 24678 1979
rect 26654 1945 26670 1979
rect 24295 1887 24528 1907
rect 26825 1887 26830 3937
rect 24295 1854 26830 1887
rect 26905 1854 26918 4311
rect 24150 1805 24187 1813
rect 21328 1784 24187 1805
rect 26899 1663 26918 1854
rect 24295 1656 26918 1663
rect 21186 1629 26918 1656
<< viali >>
rect 2669 42577 5829 42578
rect 2431 42368 5829 42577
rect 2431 42347 2752 42368
rect 2752 42347 2890 42368
rect 2890 42347 3048 42368
rect 3048 42347 3186 42368
rect 3186 42347 3344 42368
rect 3344 42347 3482 42368
rect 3482 42347 3640 42368
rect 3640 42347 3778 42368
rect 3778 42347 3936 42368
rect 3936 42347 4074 42368
rect 4074 42347 4232 42368
rect 4232 42347 4370 42368
rect 4370 42347 4528 42368
rect 4528 42347 4666 42368
rect 4666 42347 4824 42368
rect 4824 42347 4962 42368
rect 4962 42347 5120 42368
rect 5120 42347 5258 42368
rect 5258 42347 5416 42368
rect 5416 42347 5554 42368
rect 5554 42347 5829 42368
rect 2431 42272 2681 42347
rect 2431 36372 2656 42272
rect 2656 36372 2681 42272
rect 2802 41823 2840 42220
rect 2802 36424 2840 36821
rect 2431 36214 2681 36372
rect 3098 41823 3136 42220
rect 3098 36424 3136 36821
rect 3394 41823 3432 42220
rect 3394 36424 3432 36821
rect 3690 41823 3728 42220
rect 3690 36424 3728 36821
rect 3986 41823 4024 42220
rect 3986 36424 4024 36821
rect 4282 41823 4320 42220
rect 4282 36424 4320 36821
rect 4578 41823 4616 42220
rect 4578 36424 4616 36821
rect 4874 41823 4912 42220
rect 4874 36424 4912 36821
rect 5170 41823 5208 42220
rect 5170 36424 5208 36821
rect 5466 41823 5504 42220
rect 5466 36424 5504 36821
rect 5613 42272 5815 42347
rect 5613 36372 5616 42272
rect 5616 36372 5650 42272
rect 5650 36372 5815 42272
rect 2431 30314 2656 36214
rect 2656 30314 2681 36214
rect 2802 35765 2840 36162
rect 2802 30366 2840 30763
rect 2431 30245 2681 30314
rect 3098 35765 3136 36162
rect 3098 30366 3136 30763
rect 3394 35765 3432 36162
rect 3394 30366 3432 30763
rect 3690 35765 3728 36162
rect 3690 30366 3728 30763
rect 3986 35765 4024 36162
rect 3986 30366 4024 30763
rect 4282 35765 4320 36162
rect 4282 30366 4320 30763
rect 4578 35765 4616 36162
rect 4578 30366 4616 30763
rect 4874 35765 4912 36162
rect 4874 30366 4912 30763
rect 5170 35765 5208 36162
rect 5170 30366 5208 30763
rect 5466 35765 5504 36162
rect 5466 30366 5504 30763
rect 5613 36214 5815 36372
rect 5613 30314 5616 36214
rect 5616 30314 5650 36214
rect 5650 30314 5815 36214
rect 5613 30245 5815 30314
rect 2431 30218 2752 30245
rect 2752 30218 2890 30245
rect 2890 30218 3048 30245
rect 3048 30218 3186 30245
rect 3186 30218 3344 30245
rect 3344 30218 3482 30245
rect 3482 30218 3640 30245
rect 3640 30218 3778 30245
rect 3778 30218 3936 30245
rect 3936 30218 4074 30245
rect 4074 30218 4232 30245
rect 4232 30218 4370 30245
rect 4370 30218 4528 30245
rect 4528 30218 4666 30245
rect 4666 30218 4824 30245
rect 4824 30218 4962 30245
rect 4962 30218 5120 30245
rect 5120 30218 5258 30245
rect 5258 30218 5416 30245
rect 5416 30218 5554 30245
rect 5554 30218 5815 30245
rect 2431 30063 5815 30218
rect 2491 30058 5815 30063
rect 6032 31147 10883 31303
rect 6028 31137 10883 31147
rect 6028 31118 6195 31137
rect 6195 31118 8363 31137
rect 8363 31118 8521 31137
rect 8521 31118 10689 31137
rect 10689 31118 10883 31137
rect 6028 31041 6143 31118
rect 6028 30595 6099 31041
rect 6099 30595 6133 31041
rect 6133 30595 6143 31041
rect 6028 30536 6143 30595
rect 6295 30965 8263 30999
rect 6233 30730 6267 30906
rect 8291 30730 8325 30906
rect 6295 30637 8263 30671
rect 10759 31041 10874 31118
rect 8621 30965 10589 30999
rect 8559 30730 8593 30906
rect 10617 30730 10651 30906
rect 8621 30637 10589 30671
rect 10759 30595 10785 31041
rect 10785 30595 10874 31041
rect 10759 30536 10874 30595
rect 6028 30533 10882 30536
rect 6028 30499 6195 30533
rect 6195 30499 8363 30533
rect 8363 30499 8521 30533
rect 8521 30499 10689 30533
rect 10689 30499 10882 30533
rect 6028 30450 10882 30499
rect 6031 30351 10882 30450
rect 7370 28243 17591 28343
rect 7370 28209 7552 28243
rect 7552 28209 10352 28243
rect 10352 28209 10510 28243
rect 10510 28209 13310 28243
rect 13310 28230 17591 28243
rect 13310 28209 13781 28230
rect 7370 28196 13781 28209
rect 13781 28196 13815 28230
rect 13815 28196 13871 28230
rect 13871 28196 13905 28230
rect 13905 28196 13961 28230
rect 13961 28196 13995 28230
rect 13995 28196 14051 28230
rect 14051 28196 14085 28230
rect 14085 28196 14141 28230
rect 14141 28196 14175 28230
rect 14175 28196 14231 28230
rect 14231 28196 14265 28230
rect 14265 28196 14321 28230
rect 14321 28196 14355 28230
rect 14355 28196 14411 28230
rect 14411 28196 14445 28230
rect 14445 28196 14501 28230
rect 14501 28196 14535 28230
rect 14535 28196 14591 28230
rect 14591 28196 14625 28230
rect 14625 28196 14681 28230
rect 14681 28196 14715 28230
rect 14715 28196 14771 28230
rect 14771 28196 14805 28230
rect 14805 28196 15125 28230
rect 15125 28196 15159 28230
rect 15159 28196 15215 28230
rect 15215 28196 15249 28230
rect 15249 28196 15305 28230
rect 15305 28196 15339 28230
rect 15339 28196 15395 28230
rect 15395 28196 15429 28230
rect 15429 28196 15485 28230
rect 15485 28196 15519 28230
rect 15519 28196 15575 28230
rect 15575 28196 15609 28230
rect 15609 28196 15665 28230
rect 15665 28196 15699 28230
rect 15699 28196 15755 28230
rect 15755 28196 15789 28230
rect 15789 28196 15845 28230
rect 15845 28196 15879 28230
rect 15879 28196 15935 28230
rect 15935 28196 15969 28230
rect 15969 28196 16025 28230
rect 16025 28196 16059 28230
rect 16059 28196 16115 28230
rect 16115 28196 16149 28230
rect 16149 28196 16469 28230
rect 16469 28196 16503 28230
rect 16503 28196 16559 28230
rect 16559 28196 16593 28230
rect 16593 28196 16649 28230
rect 16649 28196 16683 28230
rect 16683 28196 16739 28230
rect 16739 28196 16773 28230
rect 16773 28196 16829 28230
rect 16829 28196 16863 28230
rect 16863 28196 16919 28230
rect 16919 28196 16953 28230
rect 16953 28196 17009 28230
rect 17009 28196 17043 28230
rect 17043 28196 17099 28230
rect 17099 28196 17133 28230
rect 17133 28196 17189 28230
rect 17189 28196 17223 28230
rect 17223 28196 17279 28230
rect 17279 28196 17313 28230
rect 17313 28196 17369 28230
rect 17369 28196 17403 28230
rect 17403 28196 17459 28230
rect 17459 28196 17493 28230
rect 17493 28196 17591 28230
rect 7370 28190 17591 28196
rect 7371 28147 7490 28190
rect 7371 28009 7456 28147
rect 7456 28009 7490 28147
rect 7371 27851 7490 28009
rect 7604 28059 8001 28097
rect 9903 28059 10300 28097
rect 13405 28147 17590 28190
rect 10562 28059 10959 28097
rect 12861 28059 13258 28097
rect 13405 28009 13406 28147
rect 13406 28146 17590 28147
rect 13406 28112 13680 28146
rect 13680 28112 13714 28146
rect 13714 28112 14867 28146
rect 14867 28112 14901 28146
rect 14901 28112 15024 28146
rect 15024 28112 15058 28146
rect 15058 28112 16211 28146
rect 16211 28112 16245 28146
rect 16245 28112 16368 28146
rect 16368 28112 16402 28146
rect 16402 28112 17555 28146
rect 17555 28112 17589 28146
rect 17589 28112 17590 28146
rect 13406 28080 17590 28112
rect 13406 28056 13921 28080
rect 13406 28022 13680 28056
rect 13680 28022 13714 28056
rect 13714 28050 13921 28056
rect 13921 28050 13955 28080
rect 13955 28050 14011 28080
rect 14011 28050 14045 28080
rect 14045 28050 14101 28080
rect 14101 28050 14135 28080
rect 14135 28050 14191 28080
rect 14191 28050 14225 28080
rect 14225 28050 14281 28080
rect 14281 28050 14315 28080
rect 14315 28050 14371 28080
rect 14371 28050 14405 28080
rect 14405 28050 14461 28080
rect 14461 28050 14495 28080
rect 14495 28050 14551 28080
rect 14551 28050 14585 28080
rect 14585 28050 14641 28080
rect 14641 28050 14675 28080
rect 14675 28056 15265 28080
rect 14675 28050 14867 28056
rect 13714 28022 13844 28050
rect 13406 28009 13844 28022
rect 13405 27986 13844 28009
rect 13405 27966 13829 27986
rect 13405 27932 13680 27966
rect 13680 27932 13714 27966
rect 13714 27952 13829 27966
rect 13829 27952 13844 27986
rect 14739 28022 14867 28050
rect 14867 28022 14901 28056
rect 14901 28022 15024 28056
rect 15024 28022 15058 28056
rect 15058 28050 15265 28056
rect 15265 28050 15299 28080
rect 15299 28050 15355 28080
rect 15355 28050 15389 28080
rect 15389 28050 15445 28080
rect 15445 28050 15479 28080
rect 15479 28050 15535 28080
rect 15535 28050 15569 28080
rect 15569 28050 15625 28080
rect 15625 28050 15659 28080
rect 15659 28050 15715 28080
rect 15715 28050 15749 28080
rect 15749 28050 15805 28080
rect 15805 28050 15839 28080
rect 15839 28050 15895 28080
rect 15895 28050 15929 28080
rect 15929 28050 15985 28080
rect 15985 28050 16019 28080
rect 16019 28056 16609 28080
rect 16019 28050 16211 28056
rect 15058 28022 15181 28050
rect 14739 27986 15181 28022
rect 14739 27967 15173 27986
rect 13714 27932 13844 27952
rect 13405 27896 13844 27932
rect 13405 27876 13829 27896
rect 7371 27713 7456 27851
rect 7456 27713 7490 27851
rect 7371 27555 7490 27713
rect 7604 27763 8001 27801
rect 9903 27763 10300 27801
rect 13405 27851 13680 27876
rect 10562 27763 10959 27801
rect 12861 27763 13258 27801
rect 13405 27713 13406 27851
rect 13406 27842 13680 27851
rect 13680 27842 13714 27876
rect 13714 27862 13829 27876
rect 13829 27862 13844 27896
rect 13714 27842 13844 27862
rect 13406 27806 13844 27842
rect 13406 27786 13829 27806
rect 13406 27752 13680 27786
rect 13680 27752 13714 27786
rect 13714 27772 13829 27786
rect 13829 27772 13844 27806
rect 13714 27752 13844 27772
rect 13406 27716 13844 27752
rect 13406 27713 13829 27716
rect 13405 27696 13829 27713
rect 13405 27662 13680 27696
rect 13680 27662 13714 27696
rect 13714 27682 13829 27696
rect 13829 27682 13844 27716
rect 13714 27662 13844 27682
rect 13405 27626 13844 27662
rect 13405 27606 13829 27626
rect 13405 27572 13680 27606
rect 13680 27572 13714 27606
rect 13714 27592 13829 27606
rect 13829 27592 13844 27626
rect 13714 27572 13844 27592
rect 7371 27417 7456 27555
rect 7456 27417 7490 27555
rect 7371 27259 7490 27417
rect 7604 27467 8001 27505
rect 9903 27467 10300 27505
rect 13405 27555 13844 27572
rect 10562 27467 10959 27505
rect 12861 27467 13258 27505
rect 13405 27417 13406 27555
rect 13406 27536 13844 27555
rect 13406 27516 13829 27536
rect 13406 27482 13680 27516
rect 13680 27482 13714 27516
rect 13714 27502 13829 27516
rect 13829 27502 13844 27536
rect 13714 27482 13844 27502
rect 13406 27446 13844 27482
rect 13406 27426 13829 27446
rect 13406 27417 13680 27426
rect 13405 27392 13680 27417
rect 13680 27392 13714 27426
rect 13714 27412 13829 27426
rect 13829 27412 13844 27446
rect 13714 27392 13844 27412
rect 13405 27356 13844 27392
rect 13405 27336 13829 27356
rect 13405 27302 13680 27336
rect 13680 27302 13714 27336
rect 13714 27322 13829 27336
rect 13829 27322 13844 27356
rect 13714 27302 13844 27322
rect 7371 27121 7456 27259
rect 7456 27121 7490 27259
rect 7371 26963 7490 27121
rect 7604 27171 8001 27209
rect 9903 27171 10300 27209
rect 13405 27266 13844 27302
rect 14031 27870 14037 27892
rect 14037 27870 14065 27892
rect 14031 27858 14065 27870
rect 14131 27858 14165 27892
rect 14231 27858 14265 27892
rect 14331 27870 14363 27892
rect 14363 27870 14365 27892
rect 14431 27870 14453 27892
rect 14453 27870 14465 27892
rect 14531 27870 14543 27892
rect 14543 27870 14565 27892
rect 14331 27858 14365 27870
rect 14431 27858 14465 27870
rect 14531 27858 14565 27870
rect 14031 27780 14037 27792
rect 14037 27780 14065 27792
rect 14031 27758 14065 27780
rect 14131 27758 14165 27792
rect 14231 27758 14265 27792
rect 14331 27780 14363 27792
rect 14363 27780 14365 27792
rect 14431 27780 14453 27792
rect 14453 27780 14465 27792
rect 14531 27780 14543 27792
rect 14543 27780 14565 27792
rect 14331 27758 14365 27780
rect 14431 27758 14465 27780
rect 14531 27758 14565 27780
rect 14031 27690 14037 27692
rect 14037 27690 14065 27692
rect 14031 27658 14065 27690
rect 14131 27658 14165 27692
rect 14231 27658 14265 27692
rect 14331 27690 14363 27692
rect 14363 27690 14365 27692
rect 14431 27690 14453 27692
rect 14453 27690 14465 27692
rect 14531 27690 14543 27692
rect 14543 27690 14565 27692
rect 14331 27658 14365 27690
rect 14431 27658 14465 27690
rect 14531 27658 14565 27690
rect 14031 27558 14065 27592
rect 14131 27558 14165 27592
rect 14231 27558 14265 27592
rect 14331 27558 14365 27592
rect 14431 27558 14465 27592
rect 14531 27558 14565 27592
rect 14031 27458 14065 27492
rect 14131 27458 14165 27492
rect 14231 27458 14265 27492
rect 14331 27458 14365 27492
rect 14431 27458 14465 27492
rect 14531 27458 14565 27492
rect 14031 27364 14065 27392
rect 14031 27358 14037 27364
rect 14037 27358 14065 27364
rect 14131 27358 14165 27392
rect 14231 27358 14265 27392
rect 14331 27364 14365 27392
rect 14431 27364 14465 27392
rect 14531 27364 14565 27392
rect 14331 27358 14363 27364
rect 14363 27358 14365 27364
rect 14431 27358 14453 27364
rect 14453 27358 14465 27364
rect 14531 27358 14543 27364
rect 14543 27358 14565 27364
rect 14739 27933 14753 27967
rect 14753 27966 15173 27967
rect 14753 27933 14867 27966
rect 14739 27932 14867 27933
rect 14867 27932 14901 27966
rect 14901 27932 15024 27966
rect 15024 27932 15058 27966
rect 15058 27952 15173 27966
rect 15173 27952 15181 27986
rect 16084 28022 16211 28050
rect 16211 28022 16245 28056
rect 16245 28022 16368 28056
rect 16368 28022 16402 28056
rect 16402 28050 16609 28056
rect 16609 28050 16643 28080
rect 16643 28050 16699 28080
rect 16699 28050 16733 28080
rect 16733 28050 16789 28080
rect 16789 28050 16823 28080
rect 16823 28050 16879 28080
rect 16879 28050 16913 28080
rect 16913 28050 16969 28080
rect 16969 28050 17003 28080
rect 17003 28050 17059 28080
rect 17059 28050 17093 28080
rect 17093 28050 17149 28080
rect 17149 28050 17183 28080
rect 17183 28050 17239 28080
rect 17239 28050 17273 28080
rect 17273 28050 17329 28080
rect 17329 28050 17363 28080
rect 17363 28056 17590 28080
rect 17363 28050 17555 28056
rect 16402 28022 16526 28050
rect 16084 27986 16526 28022
rect 16084 27967 16517 27986
rect 15058 27932 15181 27952
rect 14739 27896 15181 27932
rect 14739 27877 15173 27896
rect 14739 27843 14753 27877
rect 14753 27876 15173 27877
rect 14753 27843 14867 27876
rect 14739 27842 14867 27843
rect 14867 27842 14901 27876
rect 14901 27842 15024 27876
rect 15024 27842 15058 27876
rect 15058 27862 15173 27876
rect 15173 27862 15181 27896
rect 15058 27842 15181 27862
rect 14739 27825 15181 27842
rect 14762 27356 15178 27372
rect 14762 27336 15173 27356
rect 13405 27259 13829 27266
rect 10562 27171 10959 27209
rect 12861 27171 13258 27209
rect 13405 27121 13406 27259
rect 13406 27246 13829 27259
rect 13406 27212 13680 27246
rect 13680 27212 13714 27246
rect 13714 27232 13829 27246
rect 13829 27232 13844 27266
rect 13714 27212 13844 27232
rect 13406 27172 13844 27212
rect 14762 27302 14867 27336
rect 14867 27302 14901 27336
rect 14901 27302 15024 27336
rect 15024 27302 15058 27336
rect 15058 27322 15173 27336
rect 15173 27322 15178 27356
rect 15058 27302 15178 27322
rect 14762 27266 15178 27302
rect 15375 27870 15381 27892
rect 15381 27870 15409 27892
rect 15375 27858 15409 27870
rect 15475 27858 15509 27892
rect 15575 27858 15609 27892
rect 15675 27870 15707 27892
rect 15707 27870 15709 27892
rect 15775 27870 15797 27892
rect 15797 27870 15809 27892
rect 15875 27870 15887 27892
rect 15887 27870 15909 27892
rect 15675 27858 15709 27870
rect 15775 27858 15809 27870
rect 15875 27858 15909 27870
rect 15375 27780 15381 27792
rect 15381 27780 15409 27792
rect 15375 27758 15409 27780
rect 15475 27758 15509 27792
rect 15575 27758 15609 27792
rect 15675 27780 15707 27792
rect 15707 27780 15709 27792
rect 15775 27780 15797 27792
rect 15797 27780 15809 27792
rect 15875 27780 15887 27792
rect 15887 27780 15909 27792
rect 15675 27758 15709 27780
rect 15775 27758 15809 27780
rect 15875 27758 15909 27780
rect 15375 27690 15381 27692
rect 15381 27690 15409 27692
rect 15375 27658 15409 27690
rect 15475 27658 15509 27692
rect 15575 27658 15609 27692
rect 15675 27690 15707 27692
rect 15707 27690 15709 27692
rect 15775 27690 15797 27692
rect 15797 27690 15809 27692
rect 15875 27690 15887 27692
rect 15887 27690 15909 27692
rect 15675 27658 15709 27690
rect 15775 27658 15809 27690
rect 15875 27658 15909 27690
rect 15375 27558 15409 27592
rect 15475 27558 15509 27592
rect 15575 27558 15609 27592
rect 15675 27558 15709 27592
rect 15775 27558 15809 27592
rect 15875 27558 15909 27592
rect 15375 27458 15409 27492
rect 15475 27458 15509 27492
rect 15575 27458 15609 27492
rect 15675 27458 15709 27492
rect 15775 27458 15809 27492
rect 15875 27458 15909 27492
rect 15375 27364 15409 27392
rect 15375 27358 15381 27364
rect 15381 27358 15409 27364
rect 15475 27358 15509 27392
rect 15575 27358 15609 27392
rect 15675 27364 15709 27392
rect 15775 27364 15809 27392
rect 15875 27364 15909 27392
rect 15675 27358 15707 27364
rect 15707 27358 15709 27364
rect 15775 27358 15797 27364
rect 15797 27358 15809 27364
rect 15875 27358 15887 27364
rect 15887 27358 15909 27364
rect 16084 27933 16097 27967
rect 16097 27966 16517 27967
rect 16097 27933 16211 27966
rect 16084 27932 16211 27933
rect 16211 27932 16245 27966
rect 16245 27932 16368 27966
rect 16368 27932 16402 27966
rect 16402 27952 16517 27966
rect 16517 27952 16526 27986
rect 17424 28022 17555 28050
rect 17555 28022 17589 28056
rect 17589 28022 17590 28056
rect 17424 27967 17590 28022
rect 16402 27932 16526 27952
rect 16084 27896 16526 27932
rect 16084 27877 16517 27896
rect 16084 27843 16097 27877
rect 16097 27876 16517 27877
rect 16097 27843 16211 27876
rect 16084 27842 16211 27843
rect 16211 27842 16245 27876
rect 16245 27842 16368 27876
rect 16368 27842 16402 27876
rect 16402 27862 16517 27876
rect 16517 27862 16526 27896
rect 16402 27842 16526 27862
rect 16084 27814 16526 27842
rect 16092 27337 16508 27372
rect 16092 27303 16097 27337
rect 16097 27336 16508 27337
rect 16097 27303 16211 27336
rect 14762 27246 15173 27266
rect 14762 27212 14867 27246
rect 14867 27212 14901 27246
rect 14901 27212 15024 27246
rect 15024 27212 15058 27246
rect 15058 27232 15173 27246
rect 15173 27232 15178 27266
rect 15058 27212 15178 27232
rect 13406 27156 13887 27172
rect 13887 27156 13921 27172
rect 13921 27156 13977 27172
rect 13977 27156 14011 27172
rect 14011 27156 14067 27172
rect 14067 27156 14082 27172
rect 14762 27175 15178 27212
rect 16092 27302 16211 27303
rect 16211 27302 16245 27336
rect 16245 27302 16368 27336
rect 16368 27302 16402 27336
rect 16402 27302 16508 27336
rect 16092 27247 16508 27302
rect 16719 27870 16725 27892
rect 16725 27870 16753 27892
rect 16719 27858 16753 27870
rect 16819 27858 16853 27892
rect 16919 27858 16953 27892
rect 17019 27870 17051 27892
rect 17051 27870 17053 27892
rect 17119 27870 17141 27892
rect 17141 27870 17153 27892
rect 17219 27870 17231 27892
rect 17231 27870 17253 27892
rect 17019 27858 17053 27870
rect 17119 27858 17153 27870
rect 17219 27858 17253 27870
rect 16719 27780 16725 27792
rect 16725 27780 16753 27792
rect 16719 27758 16753 27780
rect 16819 27758 16853 27792
rect 16919 27758 16953 27792
rect 17019 27780 17051 27792
rect 17051 27780 17053 27792
rect 17119 27780 17141 27792
rect 17141 27780 17153 27792
rect 17219 27780 17231 27792
rect 17231 27780 17253 27792
rect 17019 27758 17053 27780
rect 17119 27758 17153 27780
rect 17219 27758 17253 27780
rect 16719 27690 16725 27692
rect 16725 27690 16753 27692
rect 16719 27658 16753 27690
rect 16819 27658 16853 27692
rect 16919 27658 16953 27692
rect 17019 27690 17051 27692
rect 17051 27690 17053 27692
rect 17119 27690 17141 27692
rect 17141 27690 17153 27692
rect 17219 27690 17231 27692
rect 17231 27690 17253 27692
rect 17019 27658 17053 27690
rect 17119 27658 17153 27690
rect 17219 27658 17253 27690
rect 16719 27558 16753 27592
rect 16819 27558 16853 27592
rect 16919 27558 16953 27592
rect 17019 27558 17053 27592
rect 17119 27558 17153 27592
rect 17219 27558 17253 27592
rect 16719 27458 16753 27492
rect 16819 27458 16853 27492
rect 16919 27458 16953 27492
rect 17019 27458 17053 27492
rect 17119 27458 17153 27492
rect 17219 27458 17253 27492
rect 16719 27364 16753 27392
rect 16719 27358 16725 27364
rect 16725 27358 16753 27364
rect 16819 27358 16853 27392
rect 16919 27358 16953 27392
rect 17019 27364 17053 27392
rect 17119 27364 17153 27392
rect 17219 27364 17253 27392
rect 17019 27358 17051 27364
rect 17051 27358 17053 27364
rect 17119 27358 17141 27364
rect 17141 27358 17153 27364
rect 17219 27358 17231 27364
rect 17231 27358 17253 27364
rect 17424 27933 17441 27967
rect 17441 27966 17590 27967
rect 17441 27933 17555 27966
rect 17424 27932 17555 27933
rect 17555 27932 17589 27966
rect 17589 27932 17590 27966
rect 17424 27877 17590 27932
rect 17424 27843 17441 27877
rect 17441 27876 17590 27877
rect 17441 27843 17555 27876
rect 17424 27842 17555 27843
rect 17555 27842 17589 27876
rect 17589 27842 17590 27876
rect 17424 27787 17590 27842
rect 17424 27753 17441 27787
rect 17441 27786 17590 27787
rect 17441 27753 17555 27786
rect 17424 27752 17555 27753
rect 17555 27752 17589 27786
rect 17589 27752 17590 27786
rect 17424 27697 17590 27752
rect 17424 27663 17441 27697
rect 17441 27696 17590 27697
rect 17441 27663 17555 27696
rect 17424 27662 17555 27663
rect 17555 27662 17589 27696
rect 17589 27662 17590 27696
rect 17424 27607 17590 27662
rect 17424 27573 17441 27607
rect 17441 27606 17590 27607
rect 17441 27573 17555 27606
rect 17424 27572 17555 27573
rect 17555 27572 17589 27606
rect 17589 27572 17590 27606
rect 17424 27517 17590 27572
rect 17424 27483 17441 27517
rect 17441 27516 17590 27517
rect 17441 27483 17555 27516
rect 17424 27482 17555 27483
rect 17555 27482 17589 27516
rect 17589 27482 17590 27516
rect 17424 27427 17590 27482
rect 17424 27393 17441 27427
rect 17441 27426 17590 27427
rect 17441 27393 17555 27426
rect 17424 27392 17555 27393
rect 17555 27392 17589 27426
rect 17589 27392 17590 27426
rect 17424 27337 17590 27392
rect 17424 27303 17441 27337
rect 17441 27336 17590 27337
rect 17441 27303 17555 27336
rect 16092 27213 16097 27247
rect 16097 27246 16508 27247
rect 16097 27213 16211 27246
rect 16092 27212 16211 27213
rect 16211 27212 16245 27246
rect 16245 27212 16368 27246
rect 16368 27212 16402 27246
rect 16402 27212 16508 27246
rect 16092 27175 16508 27212
rect 17424 27302 17555 27303
rect 17555 27302 17589 27336
rect 17589 27302 17590 27336
rect 17424 27247 17590 27302
rect 17424 27213 17441 27247
rect 17441 27246 17590 27247
rect 17441 27213 17555 27246
rect 17424 27212 17555 27213
rect 17555 27212 17589 27246
rect 17589 27212 17590 27246
rect 14550 27156 14551 27175
rect 14551 27156 14607 27175
rect 14607 27156 14641 27175
rect 14641 27156 15231 27175
rect 15231 27156 15265 27175
rect 15265 27156 15321 27175
rect 15321 27156 15355 27175
rect 15355 27156 15411 27175
rect 15411 27156 15445 27175
rect 15445 27156 15501 27175
rect 15501 27156 15535 27175
rect 15535 27156 15591 27175
rect 15591 27156 15625 27175
rect 15625 27156 15681 27175
rect 15681 27156 15715 27175
rect 15715 27156 15771 27175
rect 15771 27156 15805 27175
rect 15805 27156 15861 27175
rect 15861 27156 15895 27175
rect 15895 27156 15951 27175
rect 15951 27156 15985 27175
rect 15985 27156 16575 27175
rect 16575 27156 16609 27175
rect 16609 27156 16665 27175
rect 16665 27156 16699 27175
rect 16699 27156 16755 27175
rect 16755 27156 16764 27175
rect 17424 27179 17590 27212
rect 17195 27156 17205 27179
rect 17205 27156 17239 27179
rect 17239 27156 17295 27179
rect 17295 27156 17329 27179
rect 17329 27156 17590 27179
rect 13406 27122 13680 27156
rect 13680 27122 13714 27156
rect 13714 27122 14082 27156
rect 13406 27121 14082 27122
rect 13405 27066 14082 27121
rect 13405 27032 13680 27066
rect 13680 27032 13714 27066
rect 13714 27043 14082 27066
rect 14550 27122 14867 27156
rect 14867 27122 14901 27156
rect 14901 27122 15024 27156
rect 15024 27122 15058 27156
rect 15058 27122 16211 27156
rect 16211 27122 16245 27156
rect 16245 27122 16368 27156
rect 16368 27122 16402 27156
rect 16402 27122 16764 27156
rect 14550 27066 16764 27122
rect 14550 27043 14867 27066
rect 13714 27032 13781 27043
rect 13405 27009 13781 27032
rect 13781 27009 13815 27043
rect 13815 27009 13871 27043
rect 13871 27009 13905 27043
rect 13905 27009 13961 27043
rect 13961 27009 13995 27043
rect 13995 27009 14051 27043
rect 14051 27009 14082 27043
rect 14550 27009 14591 27043
rect 14591 27009 14625 27043
rect 14625 27009 14681 27043
rect 14681 27009 14715 27043
rect 14715 27009 14771 27043
rect 14771 27009 14805 27043
rect 14805 27032 14867 27043
rect 14867 27032 14901 27066
rect 14901 27032 15024 27066
rect 15024 27032 15058 27066
rect 15058 27043 16211 27066
rect 15058 27032 15125 27043
rect 14805 27009 15125 27032
rect 15125 27009 15159 27043
rect 15159 27009 15215 27043
rect 15215 27009 15249 27043
rect 15249 27009 15305 27043
rect 15305 27009 15339 27043
rect 15339 27009 15395 27043
rect 15395 27009 15429 27043
rect 15429 27009 15485 27043
rect 15485 27009 15519 27043
rect 15519 27009 15575 27043
rect 15575 27009 15609 27043
rect 15609 27009 15665 27043
rect 15665 27009 15699 27043
rect 15699 27009 15755 27043
rect 15755 27009 15789 27043
rect 15789 27009 15845 27043
rect 15845 27009 15879 27043
rect 15879 27009 15935 27043
rect 15935 27009 15969 27043
rect 15969 27009 16025 27043
rect 16025 27009 16059 27043
rect 16059 27009 16115 27043
rect 16115 27009 16149 27043
rect 16149 27032 16211 27043
rect 16211 27032 16245 27066
rect 16245 27032 16368 27066
rect 16368 27032 16402 27066
rect 16402 27043 16764 27066
rect 17195 27122 17555 27156
rect 17555 27122 17589 27156
rect 17589 27122 17590 27156
rect 17195 27066 17590 27122
rect 17195 27043 17555 27066
rect 16402 27032 16469 27043
rect 16149 27009 16469 27032
rect 16469 27009 16503 27043
rect 16503 27009 16559 27043
rect 16559 27009 16593 27043
rect 16593 27009 16649 27043
rect 16649 27009 16683 27043
rect 16683 27009 16739 27043
rect 16739 27009 16764 27043
rect 17195 27009 17223 27043
rect 17223 27009 17279 27043
rect 17279 27009 17313 27043
rect 17313 27009 17369 27043
rect 17369 27009 17403 27043
rect 17403 27009 17459 27043
rect 17459 27009 17493 27043
rect 17493 27032 17555 27043
rect 17555 27032 17589 27066
rect 17589 27032 17590 27066
rect 17493 27009 17590 27032
rect 7371 26825 7456 26963
rect 7456 26825 7490 26963
rect 7371 26667 7490 26825
rect 7604 26875 8001 26913
rect 9903 26875 10300 26913
rect 13405 26963 14082 27009
rect 10562 26875 10959 26913
rect 12861 26875 13258 26913
rect 13405 26825 13406 26963
rect 13406 26886 14082 26963
rect 14550 26886 16764 27009
rect 17195 26886 17590 27009
rect 13406 26852 13781 26886
rect 13781 26852 13815 26886
rect 13815 26863 13871 26886
rect 13871 26863 13905 26886
rect 13905 26863 13961 26886
rect 13961 26863 13995 26886
rect 13995 26863 14051 26886
rect 14051 26863 14082 26886
rect 13815 26852 13844 26863
rect 14550 26877 14591 26886
rect 14591 26877 14625 26886
rect 14625 26877 14681 26886
rect 14681 26877 14715 26886
rect 14715 26877 14771 26886
rect 14762 26852 14771 26877
rect 14771 26852 14805 26886
rect 14805 26852 15125 26886
rect 15125 26852 15159 26886
rect 15159 26877 15215 26886
rect 15215 26877 15249 26886
rect 15249 26877 15305 26886
rect 15305 26877 15339 26886
rect 15339 26877 15395 26886
rect 15395 26877 15429 26886
rect 15429 26877 15485 26886
rect 15485 26877 15519 26886
rect 15519 26877 15575 26886
rect 15575 26877 15609 26886
rect 15609 26877 15665 26886
rect 15665 26877 15699 26886
rect 15699 26877 15755 26886
rect 15755 26877 15789 26886
rect 15789 26877 15845 26886
rect 15845 26877 15879 26886
rect 15879 26877 15935 26886
rect 15935 26877 15969 26886
rect 15969 26877 16025 26886
rect 16025 26877 16059 26886
rect 16059 26877 16115 26886
rect 15159 26852 15178 26877
rect 16092 26852 16115 26877
rect 16115 26852 16149 26886
rect 16149 26852 16469 26886
rect 16469 26852 16503 26886
rect 16503 26877 16559 26886
rect 16559 26877 16593 26886
rect 16593 26877 16649 26886
rect 16649 26877 16683 26886
rect 16683 26877 16739 26886
rect 16739 26877 16764 26886
rect 16503 26852 16508 26877
rect 17195 26870 17223 26886
rect 17223 26870 17279 26886
rect 17279 26870 17313 26886
rect 17313 26870 17369 26886
rect 17369 26870 17403 26886
rect 17403 26870 17459 26886
rect 17424 26852 17459 26870
rect 17459 26852 17493 26886
rect 17493 26852 17590 26886
rect 13406 26825 13844 26852
rect 13405 26802 13844 26825
rect 13405 26768 13680 26802
rect 13680 26768 13714 26802
rect 13714 26768 13844 26802
rect 13405 26712 13844 26768
rect 14762 26802 15178 26852
rect 14762 26768 14867 26802
rect 14867 26768 14901 26802
rect 14901 26768 15024 26802
rect 15024 26768 15058 26802
rect 15058 26768 15178 26802
rect 7371 26529 7456 26667
rect 7456 26529 7490 26667
rect 7371 26371 7490 26529
rect 7604 26579 8001 26617
rect 9903 26579 10300 26617
rect 13405 26678 13680 26712
rect 13680 26678 13714 26712
rect 13714 26678 13844 26712
rect 14762 26712 15178 26768
rect 16092 26802 16508 26852
rect 16092 26768 16211 26802
rect 16211 26768 16245 26802
rect 16245 26768 16368 26802
rect 16368 26768 16402 26802
rect 16402 26768 16508 26802
rect 13405 26667 13844 26678
rect 10562 26579 10959 26617
rect 12861 26579 13258 26617
rect 13405 26529 13406 26667
rect 13406 26642 13844 26667
rect 13406 26622 13829 26642
rect 13406 26588 13680 26622
rect 13680 26588 13714 26622
rect 13714 26608 13829 26622
rect 13829 26608 13844 26642
rect 14762 26678 14867 26712
rect 14867 26678 14901 26712
rect 14901 26678 15024 26712
rect 15024 26678 15058 26712
rect 15058 26678 15178 26712
rect 16092 26712 16508 26768
rect 17424 26802 17590 26852
rect 17424 26768 17555 26802
rect 17555 26768 17589 26802
rect 17589 26768 17590 26802
rect 14762 26642 15178 26678
rect 13714 26588 13844 26608
rect 13406 26552 13844 26588
rect 13406 26532 13829 26552
rect 13406 26529 13680 26532
rect 13405 26498 13680 26529
rect 13680 26498 13714 26532
rect 13714 26518 13829 26532
rect 13829 26518 13844 26552
rect 13714 26498 13844 26518
rect 13405 26462 13844 26498
rect 13405 26442 13829 26462
rect 13405 26408 13680 26442
rect 13680 26408 13714 26442
rect 13714 26428 13829 26442
rect 13829 26428 13844 26462
rect 13714 26408 13844 26428
rect 7371 26233 7456 26371
rect 7456 26233 7490 26371
rect 7371 26075 7490 26233
rect 7604 26283 8001 26321
rect 9903 26283 10300 26321
rect 13405 26372 13844 26408
rect 13405 26371 13829 26372
rect 10562 26283 10959 26321
rect 12861 26283 13258 26321
rect 13405 26233 13406 26371
rect 13406 26352 13829 26371
rect 13406 26318 13680 26352
rect 13680 26318 13714 26352
rect 13714 26338 13829 26352
rect 13829 26338 13844 26372
rect 13714 26318 13844 26338
rect 13406 26282 13844 26318
rect 13406 26262 13829 26282
rect 13406 26233 13680 26262
rect 13405 26228 13680 26233
rect 13680 26228 13714 26262
rect 13714 26248 13829 26262
rect 13829 26248 13844 26282
rect 13714 26228 13844 26248
rect 13405 26192 13844 26228
rect 13405 26172 13829 26192
rect 13405 26138 13680 26172
rect 13680 26138 13714 26172
rect 13714 26158 13829 26172
rect 13829 26158 13844 26192
rect 13714 26138 13844 26158
rect 13405 26102 13844 26138
rect 7371 25937 7456 26075
rect 7456 25937 7490 26075
rect 7371 25779 7490 25937
rect 7604 25987 8001 26025
rect 9903 25987 10300 26025
rect 13405 26082 13829 26102
rect 13405 26075 13680 26082
rect 10562 25987 10959 26025
rect 12861 25987 13258 26025
rect 13405 25937 13406 26075
rect 13406 26048 13680 26075
rect 13680 26048 13714 26082
rect 13714 26068 13829 26082
rect 13829 26068 13844 26102
rect 13714 26048 13844 26068
rect 13406 26012 13844 26048
rect 13406 25992 13829 26012
rect 13406 25958 13680 25992
rect 13680 25958 13714 25992
rect 13714 25978 13829 25992
rect 13829 25978 13844 26012
rect 13714 25958 13844 25978
rect 13406 25937 13844 25958
rect 13405 25922 13844 25937
rect 14031 26526 14037 26548
rect 14037 26526 14065 26548
rect 14031 26514 14065 26526
rect 14131 26514 14165 26548
rect 14231 26514 14265 26548
rect 14331 26526 14363 26548
rect 14363 26526 14365 26548
rect 14431 26526 14453 26548
rect 14453 26526 14465 26548
rect 14531 26526 14543 26548
rect 14543 26526 14565 26548
rect 14331 26514 14365 26526
rect 14431 26514 14465 26526
rect 14531 26514 14565 26526
rect 14031 26436 14037 26448
rect 14037 26436 14065 26448
rect 14031 26414 14065 26436
rect 14131 26414 14165 26448
rect 14231 26414 14265 26448
rect 14331 26436 14363 26448
rect 14363 26436 14365 26448
rect 14431 26436 14453 26448
rect 14453 26436 14465 26448
rect 14531 26436 14543 26448
rect 14543 26436 14565 26448
rect 14331 26414 14365 26436
rect 14431 26414 14465 26436
rect 14531 26414 14565 26436
rect 14031 26346 14037 26348
rect 14037 26346 14065 26348
rect 14031 26314 14065 26346
rect 14131 26314 14165 26348
rect 14231 26314 14265 26348
rect 14331 26346 14363 26348
rect 14363 26346 14365 26348
rect 14431 26346 14453 26348
rect 14453 26346 14465 26348
rect 14531 26346 14543 26348
rect 14543 26346 14565 26348
rect 14331 26314 14365 26346
rect 14431 26314 14465 26346
rect 14531 26314 14565 26346
rect 14031 26214 14065 26248
rect 14131 26214 14165 26248
rect 14231 26214 14265 26248
rect 14331 26214 14365 26248
rect 14431 26214 14465 26248
rect 14531 26214 14565 26248
rect 14031 26114 14065 26148
rect 14131 26114 14165 26148
rect 14231 26114 14265 26148
rect 14331 26114 14365 26148
rect 14431 26114 14465 26148
rect 14531 26114 14565 26148
rect 14031 26020 14065 26048
rect 14031 26014 14037 26020
rect 14037 26014 14065 26020
rect 14131 26014 14165 26048
rect 14231 26014 14265 26048
rect 14331 26020 14365 26048
rect 14431 26020 14465 26048
rect 14531 26020 14565 26048
rect 14331 26014 14363 26020
rect 14363 26014 14365 26020
rect 14431 26014 14453 26020
rect 14453 26014 14465 26020
rect 14531 26014 14543 26020
rect 14543 26014 14565 26020
rect 14762 26622 15173 26642
rect 14762 26588 14867 26622
rect 14867 26588 14901 26622
rect 14901 26588 15024 26622
rect 15024 26588 15058 26622
rect 15058 26608 15173 26622
rect 15173 26608 15178 26642
rect 16092 26678 16211 26712
rect 16211 26678 16245 26712
rect 16245 26678 16368 26712
rect 16368 26678 16402 26712
rect 16402 26678 16508 26712
rect 17424 26712 17590 26768
rect 16092 26623 16508 26678
rect 15058 26588 15178 26608
rect 14762 26552 15178 26588
rect 14762 26532 15173 26552
rect 14762 26498 14867 26532
rect 14867 26498 14901 26532
rect 14901 26498 15024 26532
rect 15024 26498 15058 26532
rect 15058 26518 15173 26532
rect 15173 26518 15178 26552
rect 15058 26498 15178 26518
rect 14762 26462 15178 26498
rect 14762 26442 15173 26462
rect 14762 26408 14867 26442
rect 14867 26408 14901 26442
rect 14901 26408 15024 26442
rect 15024 26408 15058 26442
rect 15058 26428 15173 26442
rect 15173 26428 15178 26462
rect 15058 26408 15178 26428
rect 14762 26372 15178 26408
rect 14762 26352 15173 26372
rect 14762 26318 14867 26352
rect 14867 26318 14901 26352
rect 14901 26318 15024 26352
rect 15024 26318 15058 26352
rect 15058 26338 15173 26352
rect 15173 26338 15178 26372
rect 15058 26318 15178 26338
rect 14762 26282 15178 26318
rect 14762 26262 15173 26282
rect 14762 26228 14867 26262
rect 14867 26228 14901 26262
rect 14901 26228 15024 26262
rect 15024 26228 15058 26262
rect 15058 26248 15173 26262
rect 15173 26248 15178 26282
rect 15058 26228 15178 26248
rect 14762 26192 15178 26228
rect 14762 26172 15173 26192
rect 14762 26138 14867 26172
rect 14867 26138 14901 26172
rect 14901 26138 15024 26172
rect 15024 26138 15058 26172
rect 15058 26158 15173 26172
rect 15173 26158 15178 26192
rect 15058 26138 15178 26158
rect 14762 26102 15178 26138
rect 14762 26082 15173 26102
rect 14762 26048 14867 26082
rect 14867 26048 14901 26082
rect 14901 26048 15024 26082
rect 15024 26048 15058 26082
rect 15058 26068 15173 26082
rect 15173 26068 15178 26102
rect 15058 26048 15178 26068
rect 14762 26012 15178 26048
rect 14762 25992 15173 26012
rect 13405 25902 13829 25922
rect 13405 25868 13680 25902
rect 13680 25868 13714 25902
rect 13714 25888 13829 25902
rect 13829 25888 13844 25922
rect 13714 25868 13844 25888
rect 13405 25826 13844 25868
rect 14762 25958 14867 25992
rect 14867 25958 14901 25992
rect 14901 25958 15024 25992
rect 15024 25958 15058 25992
rect 15058 25978 15173 25992
rect 15173 25978 15178 26012
rect 15058 25958 15178 25978
rect 14762 25922 15178 25958
rect 15375 26526 15381 26548
rect 15381 26526 15409 26548
rect 15375 26514 15409 26526
rect 15475 26514 15509 26548
rect 15575 26514 15609 26548
rect 15675 26526 15707 26548
rect 15707 26526 15709 26548
rect 15775 26526 15797 26548
rect 15797 26526 15809 26548
rect 15875 26526 15887 26548
rect 15887 26526 15909 26548
rect 15675 26514 15709 26526
rect 15775 26514 15809 26526
rect 15875 26514 15909 26526
rect 15375 26436 15381 26448
rect 15381 26436 15409 26448
rect 15375 26414 15409 26436
rect 15475 26414 15509 26448
rect 15575 26414 15609 26448
rect 15675 26436 15707 26448
rect 15707 26436 15709 26448
rect 15775 26436 15797 26448
rect 15797 26436 15809 26448
rect 15875 26436 15887 26448
rect 15887 26436 15909 26448
rect 15675 26414 15709 26436
rect 15775 26414 15809 26436
rect 15875 26414 15909 26436
rect 15375 26346 15381 26348
rect 15381 26346 15409 26348
rect 15375 26314 15409 26346
rect 15475 26314 15509 26348
rect 15575 26314 15609 26348
rect 15675 26346 15707 26348
rect 15707 26346 15709 26348
rect 15775 26346 15797 26348
rect 15797 26346 15809 26348
rect 15875 26346 15887 26348
rect 15887 26346 15909 26348
rect 15675 26314 15709 26346
rect 15775 26314 15809 26346
rect 15875 26314 15909 26346
rect 15375 26214 15409 26248
rect 15475 26214 15509 26248
rect 15575 26214 15609 26248
rect 15675 26214 15709 26248
rect 15775 26214 15809 26248
rect 15875 26214 15909 26248
rect 15375 26114 15409 26148
rect 15475 26114 15509 26148
rect 15575 26114 15609 26148
rect 15675 26114 15709 26148
rect 15775 26114 15809 26148
rect 15875 26114 15909 26148
rect 15375 26020 15409 26048
rect 15375 26014 15381 26020
rect 15381 26014 15409 26020
rect 15475 26014 15509 26048
rect 15575 26014 15609 26048
rect 15675 26020 15709 26048
rect 15775 26020 15809 26048
rect 15875 26020 15909 26048
rect 15675 26014 15707 26020
rect 15707 26014 15709 26020
rect 15775 26014 15797 26020
rect 15797 26014 15809 26020
rect 15875 26014 15887 26020
rect 15887 26014 15909 26020
rect 16092 26589 16097 26623
rect 16097 26622 16508 26623
rect 16097 26589 16211 26622
rect 16092 26588 16211 26589
rect 16211 26588 16245 26622
rect 16245 26588 16368 26622
rect 16368 26588 16402 26622
rect 16402 26588 16508 26622
rect 17424 26678 17555 26712
rect 17555 26678 17589 26712
rect 17589 26678 17590 26712
rect 17424 26623 17590 26678
rect 16092 26533 16508 26588
rect 16092 26499 16097 26533
rect 16097 26532 16508 26533
rect 16097 26499 16211 26532
rect 16092 26498 16211 26499
rect 16211 26498 16245 26532
rect 16245 26498 16368 26532
rect 16368 26498 16402 26532
rect 16402 26498 16508 26532
rect 16092 26443 16508 26498
rect 16092 26409 16097 26443
rect 16097 26442 16508 26443
rect 16097 26409 16211 26442
rect 16092 26408 16211 26409
rect 16211 26408 16245 26442
rect 16245 26408 16368 26442
rect 16368 26408 16402 26442
rect 16402 26408 16508 26442
rect 16092 26353 16508 26408
rect 16092 26319 16097 26353
rect 16097 26352 16508 26353
rect 16097 26319 16211 26352
rect 16092 26318 16211 26319
rect 16211 26318 16245 26352
rect 16245 26318 16368 26352
rect 16368 26318 16402 26352
rect 16402 26318 16508 26352
rect 16092 26263 16508 26318
rect 16092 26229 16097 26263
rect 16097 26262 16508 26263
rect 16097 26229 16211 26262
rect 16092 26228 16211 26229
rect 16211 26228 16245 26262
rect 16245 26228 16368 26262
rect 16368 26228 16402 26262
rect 16402 26228 16508 26262
rect 16092 26173 16508 26228
rect 16092 26139 16097 26173
rect 16097 26172 16508 26173
rect 16097 26139 16211 26172
rect 16092 26138 16211 26139
rect 16211 26138 16245 26172
rect 16245 26138 16368 26172
rect 16368 26138 16402 26172
rect 16402 26138 16508 26172
rect 16092 26083 16508 26138
rect 16092 26049 16097 26083
rect 16097 26082 16508 26083
rect 16097 26049 16211 26082
rect 16092 26048 16211 26049
rect 16211 26048 16245 26082
rect 16245 26048 16368 26082
rect 16368 26048 16402 26082
rect 16402 26048 16508 26082
rect 16092 25993 16508 26048
rect 16092 25959 16097 25993
rect 16097 25992 16508 25993
rect 16097 25959 16211 25992
rect 14762 25902 15173 25922
rect 14762 25868 14867 25902
rect 14867 25868 14901 25902
rect 14901 25868 15024 25902
rect 15024 25868 15058 25902
rect 15058 25888 15173 25902
rect 15173 25888 15178 25922
rect 15058 25868 15178 25888
rect 13405 25812 13887 25826
rect 13887 25812 13921 25826
rect 13921 25812 13977 25826
rect 13977 25812 14011 25826
rect 14011 25812 14067 25826
rect 14067 25812 14082 25826
rect 14762 25826 15178 25868
rect 16092 25958 16211 25959
rect 16211 25958 16245 25992
rect 16245 25958 16368 25992
rect 16368 25958 16402 25992
rect 16402 25958 16508 25992
rect 16092 25903 16508 25958
rect 16719 26526 16725 26548
rect 16725 26526 16753 26548
rect 16719 26514 16753 26526
rect 16819 26514 16853 26548
rect 16919 26514 16953 26548
rect 17019 26526 17051 26548
rect 17051 26526 17053 26548
rect 17119 26526 17141 26548
rect 17141 26526 17153 26548
rect 17219 26526 17231 26548
rect 17231 26526 17253 26548
rect 17019 26514 17053 26526
rect 17119 26514 17153 26526
rect 17219 26514 17253 26526
rect 16719 26436 16725 26448
rect 16725 26436 16753 26448
rect 16719 26414 16753 26436
rect 16819 26414 16853 26448
rect 16919 26414 16953 26448
rect 17019 26436 17051 26448
rect 17051 26436 17053 26448
rect 17119 26436 17141 26448
rect 17141 26436 17153 26448
rect 17219 26436 17231 26448
rect 17231 26436 17253 26448
rect 17019 26414 17053 26436
rect 17119 26414 17153 26436
rect 17219 26414 17253 26436
rect 16719 26346 16725 26348
rect 16725 26346 16753 26348
rect 16719 26314 16753 26346
rect 16819 26314 16853 26348
rect 16919 26314 16953 26348
rect 17019 26346 17051 26348
rect 17051 26346 17053 26348
rect 17119 26346 17141 26348
rect 17141 26346 17153 26348
rect 17219 26346 17231 26348
rect 17231 26346 17253 26348
rect 17019 26314 17053 26346
rect 17119 26314 17153 26346
rect 17219 26314 17253 26346
rect 16719 26214 16753 26248
rect 16819 26214 16853 26248
rect 16919 26214 16953 26248
rect 17019 26214 17053 26248
rect 17119 26214 17153 26248
rect 17219 26214 17253 26248
rect 16719 26114 16753 26148
rect 16819 26114 16853 26148
rect 16919 26114 16953 26148
rect 17019 26114 17053 26148
rect 17119 26114 17153 26148
rect 17219 26114 17253 26148
rect 16719 26020 16753 26048
rect 16719 26014 16725 26020
rect 16725 26014 16753 26020
rect 16819 26014 16853 26048
rect 16919 26014 16953 26048
rect 17019 26020 17053 26048
rect 17119 26020 17153 26048
rect 17219 26020 17253 26048
rect 17019 26014 17051 26020
rect 17051 26014 17053 26020
rect 17119 26014 17141 26020
rect 17141 26014 17153 26020
rect 17219 26014 17231 26020
rect 17231 26014 17253 26020
rect 17424 26589 17441 26623
rect 17441 26622 17590 26623
rect 17441 26589 17555 26622
rect 17424 26588 17555 26589
rect 17555 26588 17589 26622
rect 17589 26588 17590 26622
rect 17424 26533 17590 26588
rect 17424 26499 17441 26533
rect 17441 26532 17590 26533
rect 17441 26499 17555 26532
rect 17424 26498 17555 26499
rect 17555 26498 17589 26532
rect 17589 26498 17590 26532
rect 17424 26443 17590 26498
rect 17424 26409 17441 26443
rect 17441 26442 17590 26443
rect 17441 26409 17555 26442
rect 17424 26408 17555 26409
rect 17555 26408 17589 26442
rect 17589 26408 17590 26442
rect 17424 26353 17590 26408
rect 17424 26319 17441 26353
rect 17441 26352 17590 26353
rect 17441 26319 17555 26352
rect 17424 26318 17555 26319
rect 17555 26318 17589 26352
rect 17589 26318 17590 26352
rect 17424 26263 17590 26318
rect 17424 26229 17441 26263
rect 17441 26262 17590 26263
rect 17441 26229 17555 26262
rect 17424 26228 17555 26229
rect 17555 26228 17589 26262
rect 17589 26228 17590 26262
rect 17424 26173 17590 26228
rect 17424 26139 17441 26173
rect 17441 26172 17590 26173
rect 17441 26139 17555 26172
rect 17424 26138 17555 26139
rect 17555 26138 17589 26172
rect 17589 26138 17590 26172
rect 17424 26083 17590 26138
rect 17424 26049 17441 26083
rect 17441 26082 17590 26083
rect 17441 26049 17555 26082
rect 17424 26048 17555 26049
rect 17555 26048 17589 26082
rect 17589 26048 17590 26082
rect 17424 25993 17590 26048
rect 17424 25959 17441 25993
rect 17441 25992 17590 25993
rect 17441 25959 17555 25992
rect 16092 25869 16097 25903
rect 16097 25902 16508 25903
rect 16097 25869 16211 25902
rect 16092 25868 16211 25869
rect 16211 25868 16245 25902
rect 16245 25868 16368 25902
rect 16368 25868 16402 25902
rect 16402 25868 16508 25902
rect 16092 25826 16508 25868
rect 17424 25958 17555 25959
rect 17555 25958 17589 25992
rect 17589 25958 17590 25992
rect 17424 25903 17590 25958
rect 17424 25869 17441 25903
rect 17441 25902 17590 25903
rect 17441 25869 17555 25902
rect 17424 25868 17555 25869
rect 17555 25868 17589 25902
rect 17589 25868 17590 25902
rect 14581 25812 14607 25826
rect 14607 25812 14641 25826
rect 14641 25812 15231 25826
rect 15231 25812 15265 25826
rect 15265 25812 15321 25826
rect 15321 25812 15355 25826
rect 15355 25812 15411 25826
rect 15411 25812 15445 25826
rect 15445 25812 15501 25826
rect 15501 25812 15535 25826
rect 15535 25812 15591 25826
rect 15591 25812 15625 25826
rect 15625 25812 15681 25826
rect 15681 25812 15715 25826
rect 15715 25812 15771 25826
rect 15771 25812 15805 25826
rect 15805 25812 15861 25826
rect 15861 25812 15895 25826
rect 15895 25812 15951 25826
rect 15951 25812 15985 25826
rect 15985 25812 16575 25826
rect 16575 25812 16609 25826
rect 16609 25812 16665 25826
rect 16665 25812 16699 25826
rect 16699 25812 16753 25826
rect 17424 25845 17590 25868
rect 17210 25812 17239 25845
rect 17239 25812 17295 25845
rect 17295 25812 17329 25845
rect 17329 25812 17590 25845
rect 7371 25641 7456 25779
rect 7456 25641 7490 25779
rect 7371 25483 7490 25641
rect 7604 25691 8001 25729
rect 9903 25691 10300 25729
rect 13405 25779 13680 25812
rect 10562 25691 10959 25729
rect 12861 25691 13258 25729
rect 13405 25641 13406 25779
rect 13406 25778 13680 25779
rect 13680 25778 13714 25812
rect 13714 25778 14082 25812
rect 13406 25722 14082 25778
rect 13406 25688 13680 25722
rect 13680 25688 13714 25722
rect 13714 25699 14082 25722
rect 14581 25778 14867 25812
rect 14867 25778 14901 25812
rect 14901 25778 15024 25812
rect 15024 25778 15058 25812
rect 15058 25778 16211 25812
rect 16211 25778 16245 25812
rect 16245 25778 16368 25812
rect 16368 25778 16402 25812
rect 16402 25778 16753 25812
rect 14581 25722 16753 25778
rect 14581 25699 14867 25722
rect 13714 25688 13781 25699
rect 13406 25665 13781 25688
rect 13781 25665 13815 25699
rect 13815 25665 13871 25699
rect 13871 25665 13905 25699
rect 13905 25665 13961 25699
rect 13961 25665 13995 25699
rect 13995 25665 14051 25699
rect 14051 25665 14082 25699
rect 14581 25665 14591 25699
rect 14591 25665 14625 25699
rect 14625 25665 14681 25699
rect 14681 25665 14715 25699
rect 14715 25665 14771 25699
rect 14771 25665 14805 25699
rect 14805 25688 14867 25699
rect 14867 25688 14901 25722
rect 14901 25688 15024 25722
rect 15024 25688 15058 25722
rect 15058 25699 16211 25722
rect 15058 25688 15125 25699
rect 14805 25665 15125 25688
rect 15125 25665 15159 25699
rect 15159 25665 15215 25699
rect 15215 25665 15249 25699
rect 15249 25665 15305 25699
rect 15305 25665 15339 25699
rect 15339 25665 15395 25699
rect 15395 25665 15429 25699
rect 15429 25665 15485 25699
rect 15485 25665 15519 25699
rect 15519 25665 15575 25699
rect 15575 25665 15609 25699
rect 15609 25665 15665 25699
rect 15665 25665 15699 25699
rect 15699 25665 15755 25699
rect 15755 25665 15789 25699
rect 15789 25665 15845 25699
rect 15845 25665 15879 25699
rect 15879 25665 15935 25699
rect 15935 25665 15969 25699
rect 15969 25665 16025 25699
rect 16025 25665 16059 25699
rect 16059 25665 16115 25699
rect 16115 25665 16149 25699
rect 16149 25688 16211 25699
rect 16211 25688 16245 25722
rect 16245 25688 16368 25722
rect 16368 25688 16402 25722
rect 16402 25699 16753 25722
rect 17210 25778 17555 25812
rect 17555 25778 17589 25812
rect 17589 25778 17590 25812
rect 17210 25722 17590 25778
rect 17210 25699 17555 25722
rect 16402 25688 16469 25699
rect 16149 25665 16469 25688
rect 16469 25665 16503 25699
rect 16503 25665 16559 25699
rect 16559 25665 16593 25699
rect 16593 25665 16649 25699
rect 16649 25665 16683 25699
rect 16683 25665 16739 25699
rect 16739 25665 16753 25699
rect 17210 25665 17223 25699
rect 17223 25665 17279 25699
rect 17279 25665 17313 25699
rect 17313 25665 17369 25699
rect 17369 25665 17403 25699
rect 17403 25665 17459 25699
rect 17459 25665 17493 25699
rect 17493 25688 17555 25699
rect 17555 25688 17589 25722
rect 17589 25688 17590 25722
rect 17493 25665 17590 25688
rect 13406 25641 14082 25665
rect 13405 25542 14082 25641
rect 14581 25542 16753 25665
rect 17210 25542 17590 25665
rect 13405 25508 13781 25542
rect 13781 25508 13815 25542
rect 13815 25517 13871 25542
rect 13871 25517 13905 25542
rect 13905 25517 13961 25542
rect 13961 25517 13995 25542
rect 13995 25517 14051 25542
rect 14051 25517 14082 25542
rect 13815 25508 13844 25517
rect 14581 25520 14591 25542
rect 14591 25520 14625 25542
rect 14625 25520 14681 25542
rect 14681 25520 14715 25542
rect 14715 25520 14771 25542
rect 14762 25508 14771 25520
rect 14771 25508 14805 25542
rect 14805 25508 15125 25542
rect 15125 25508 15159 25542
rect 15159 25520 15215 25542
rect 15215 25520 15249 25542
rect 15249 25520 15305 25542
rect 15305 25520 15339 25542
rect 15339 25520 15395 25542
rect 15395 25520 15429 25542
rect 15429 25520 15485 25542
rect 15485 25520 15519 25542
rect 15519 25520 15575 25542
rect 15575 25520 15609 25542
rect 15609 25520 15665 25542
rect 15665 25520 15699 25542
rect 15699 25520 15755 25542
rect 15755 25520 15789 25542
rect 15789 25520 15845 25542
rect 15845 25520 15879 25542
rect 15879 25520 15935 25542
rect 15935 25520 15969 25542
rect 15969 25520 16025 25542
rect 16025 25520 16059 25542
rect 16059 25520 16115 25542
rect 15159 25508 15178 25520
rect 16092 25508 16115 25520
rect 16115 25508 16149 25542
rect 16149 25508 16469 25542
rect 16469 25508 16503 25542
rect 16503 25520 16559 25542
rect 16559 25520 16593 25542
rect 16593 25520 16649 25542
rect 16649 25520 16683 25542
rect 16683 25520 16739 25542
rect 16739 25520 16753 25542
rect 16503 25508 16508 25520
rect 17210 25508 17223 25542
rect 17223 25508 17279 25542
rect 17279 25508 17313 25542
rect 17313 25508 17369 25542
rect 17369 25508 17403 25542
rect 17403 25508 17459 25542
rect 17459 25508 17493 25542
rect 17493 25508 17590 25542
rect 7371 25345 7456 25483
rect 7456 25345 7490 25483
rect 7371 25187 7490 25345
rect 7604 25395 8001 25433
rect 9903 25395 10300 25433
rect 13405 25483 13844 25508
rect 10562 25395 10959 25433
rect 12861 25395 13258 25433
rect 13405 25345 13406 25483
rect 13406 25458 13844 25483
rect 13406 25424 13680 25458
rect 13680 25424 13714 25458
rect 13714 25424 13844 25458
rect 13406 25368 13844 25424
rect 14762 25458 15178 25508
rect 14762 25424 14867 25458
rect 14867 25424 14901 25458
rect 14901 25424 15024 25458
rect 15024 25424 15058 25458
rect 15058 25424 15178 25458
rect 13406 25345 13680 25368
rect 13405 25334 13680 25345
rect 13680 25334 13714 25368
rect 13714 25334 13844 25368
rect 14762 25368 15178 25424
rect 16092 25458 16508 25508
rect 17210 25501 17590 25508
rect 16092 25424 16211 25458
rect 16211 25424 16245 25458
rect 16245 25424 16368 25458
rect 16368 25424 16402 25458
rect 16402 25424 16508 25458
rect 13405 25298 13844 25334
rect 13405 25278 13829 25298
rect 13405 25244 13680 25278
rect 13680 25244 13714 25278
rect 13714 25264 13829 25278
rect 13829 25264 13844 25298
rect 14762 25334 14867 25368
rect 14867 25334 14901 25368
rect 14901 25334 15024 25368
rect 15024 25334 15058 25368
rect 15058 25334 15178 25368
rect 16092 25368 16508 25424
rect 17424 25458 17590 25501
rect 17424 25424 17555 25458
rect 17555 25424 17589 25458
rect 17589 25424 17590 25458
rect 14762 25298 15178 25334
rect 13714 25244 13844 25264
rect 7371 25049 7456 25187
rect 7456 25049 7490 25187
rect 7371 24891 7490 25049
rect 7604 25099 8001 25137
rect 9903 25099 10300 25137
rect 13405 25208 13844 25244
rect 13405 25188 13829 25208
rect 13405 25187 13680 25188
rect 10562 25099 10959 25137
rect 12861 25099 13258 25137
rect 13405 25049 13406 25187
rect 13406 25154 13680 25187
rect 13680 25154 13714 25188
rect 13714 25174 13829 25188
rect 13829 25174 13844 25208
rect 13714 25154 13844 25174
rect 13406 25118 13844 25154
rect 13406 25098 13829 25118
rect 13406 25064 13680 25098
rect 13680 25064 13714 25098
rect 13714 25084 13829 25098
rect 13829 25084 13844 25118
rect 13714 25064 13844 25084
rect 13406 25049 13844 25064
rect 13405 25028 13844 25049
rect 13405 25008 13829 25028
rect 13405 24974 13680 25008
rect 13680 24974 13714 25008
rect 13714 24994 13829 25008
rect 13829 24994 13844 25028
rect 13714 24974 13844 24994
rect 13405 24938 13844 24974
rect 13405 24918 13829 24938
rect 7371 24753 7456 24891
rect 7456 24753 7490 24891
rect 5742 24614 5981 24621
rect 7371 24614 7490 24753
rect 7604 24803 8001 24841
rect 9903 24803 10300 24841
rect 13405 24891 13680 24918
rect 10562 24803 10959 24841
rect 12861 24803 13258 24841
rect 13405 24753 13406 24891
rect 13406 24884 13680 24891
rect 13680 24884 13714 24918
rect 13714 24904 13829 24918
rect 13829 24904 13844 24938
rect 13714 24884 13844 24904
rect 13406 24848 13844 24884
rect 13406 24828 13829 24848
rect 13406 24794 13680 24828
rect 13680 24794 13714 24828
rect 13714 24814 13829 24828
rect 13829 24814 13844 24848
rect 13714 24794 13844 24814
rect 13406 24758 13844 24794
rect 13406 24753 13829 24758
rect 13405 24738 13829 24753
rect 13405 24704 13680 24738
rect 13680 24704 13714 24738
rect 13714 24724 13829 24738
rect 13829 24724 13844 24758
rect 13714 24704 13844 24724
rect 13405 24668 13844 24704
rect 13405 24648 13829 24668
rect 13405 24614 13680 24648
rect 13680 24614 13714 24648
rect 13714 24634 13829 24648
rect 13829 24634 13844 24668
rect 13714 24614 13844 24634
rect 5742 24602 11232 24614
rect 13405 24602 13844 24614
rect 5742 24578 13844 24602
rect 14031 25182 14037 25204
rect 14037 25182 14065 25204
rect 14031 25170 14065 25182
rect 14131 25170 14165 25204
rect 14231 25170 14265 25204
rect 14331 25182 14363 25204
rect 14363 25182 14365 25204
rect 14431 25182 14453 25204
rect 14453 25182 14465 25204
rect 14531 25182 14543 25204
rect 14543 25182 14565 25204
rect 14331 25170 14365 25182
rect 14431 25170 14465 25182
rect 14531 25170 14565 25182
rect 14031 25092 14037 25104
rect 14037 25092 14065 25104
rect 14031 25070 14065 25092
rect 14131 25070 14165 25104
rect 14231 25070 14265 25104
rect 14331 25092 14363 25104
rect 14363 25092 14365 25104
rect 14431 25092 14453 25104
rect 14453 25092 14465 25104
rect 14531 25092 14543 25104
rect 14543 25092 14565 25104
rect 14331 25070 14365 25092
rect 14431 25070 14465 25092
rect 14531 25070 14565 25092
rect 14031 25002 14037 25004
rect 14037 25002 14065 25004
rect 14031 24970 14065 25002
rect 14131 24970 14165 25004
rect 14231 24970 14265 25004
rect 14331 25002 14363 25004
rect 14363 25002 14365 25004
rect 14431 25002 14453 25004
rect 14453 25002 14465 25004
rect 14531 25002 14543 25004
rect 14543 25002 14565 25004
rect 14331 24970 14365 25002
rect 14431 24970 14465 25002
rect 14531 24970 14565 25002
rect 14031 24870 14065 24904
rect 14131 24870 14165 24904
rect 14231 24870 14265 24904
rect 14331 24870 14365 24904
rect 14431 24870 14465 24904
rect 14531 24870 14565 24904
rect 14031 24770 14065 24804
rect 14131 24770 14165 24804
rect 14231 24770 14265 24804
rect 14331 24770 14365 24804
rect 14431 24770 14465 24804
rect 14531 24770 14565 24804
rect 14031 24676 14065 24704
rect 14031 24670 14037 24676
rect 14037 24670 14065 24676
rect 14131 24670 14165 24704
rect 14231 24670 14265 24704
rect 14331 24676 14365 24704
rect 14431 24676 14465 24704
rect 14531 24676 14565 24704
rect 14331 24670 14363 24676
rect 14363 24670 14365 24676
rect 14431 24670 14453 24676
rect 14453 24670 14465 24676
rect 14531 24670 14543 24676
rect 14543 24670 14565 24676
rect 14762 25278 15173 25298
rect 14762 25244 14867 25278
rect 14867 25244 14901 25278
rect 14901 25244 15024 25278
rect 15024 25244 15058 25278
rect 15058 25264 15173 25278
rect 15173 25264 15178 25298
rect 16092 25334 16211 25368
rect 16211 25334 16245 25368
rect 16245 25334 16368 25368
rect 16368 25334 16402 25368
rect 16402 25334 16508 25368
rect 17424 25368 17590 25424
rect 16092 25279 16508 25334
rect 15058 25244 15178 25264
rect 14762 25208 15178 25244
rect 14762 25188 15173 25208
rect 14762 25154 14867 25188
rect 14867 25154 14901 25188
rect 14901 25154 15024 25188
rect 15024 25154 15058 25188
rect 15058 25174 15173 25188
rect 15173 25174 15178 25208
rect 15058 25154 15178 25174
rect 14762 25118 15178 25154
rect 14762 25105 15173 25118
rect 15173 25105 15178 25118
rect 14743 24705 14753 24716
rect 14753 24705 14867 24716
rect 14743 24704 14867 24705
rect 14867 24704 14901 24716
rect 14901 24704 15024 24716
rect 15024 24704 15058 24716
rect 15058 24704 15185 24716
rect 14743 24668 15185 24704
rect 14743 24649 15173 24668
rect 14743 24615 14753 24649
rect 14753 24648 15173 24649
rect 14753 24615 14867 24648
rect 5742 24558 13829 24578
rect 5742 24524 13680 24558
rect 13680 24524 13714 24558
rect 13714 24544 13829 24558
rect 13829 24544 13844 24578
rect 13714 24524 13844 24544
rect 5742 24496 13844 24524
rect 14743 24614 14867 24615
rect 14867 24614 14901 24648
rect 14901 24614 15024 24648
rect 15024 24614 15058 24648
rect 15058 24634 15173 24648
rect 15173 24634 15185 24668
rect 15058 24614 15185 24634
rect 14743 24578 15185 24614
rect 15375 25182 15381 25204
rect 15381 25182 15409 25204
rect 15375 25170 15409 25182
rect 15475 25170 15509 25204
rect 15575 25170 15609 25204
rect 15675 25182 15707 25204
rect 15707 25182 15709 25204
rect 15775 25182 15797 25204
rect 15797 25182 15809 25204
rect 15875 25182 15887 25204
rect 15887 25182 15909 25204
rect 15675 25170 15709 25182
rect 15775 25170 15809 25182
rect 15875 25170 15909 25182
rect 15375 25092 15381 25104
rect 15381 25092 15409 25104
rect 15375 25070 15409 25092
rect 15475 25070 15509 25104
rect 15575 25070 15609 25104
rect 15675 25092 15707 25104
rect 15707 25092 15709 25104
rect 15775 25092 15797 25104
rect 15797 25092 15809 25104
rect 15875 25092 15887 25104
rect 15887 25092 15909 25104
rect 15675 25070 15709 25092
rect 15775 25070 15809 25092
rect 15875 25070 15909 25092
rect 15375 25002 15381 25004
rect 15381 25002 15409 25004
rect 15375 24970 15409 25002
rect 15475 24970 15509 25004
rect 15575 24970 15609 25004
rect 15675 25002 15707 25004
rect 15707 25002 15709 25004
rect 15775 25002 15797 25004
rect 15797 25002 15809 25004
rect 15875 25002 15887 25004
rect 15887 25002 15909 25004
rect 15675 24970 15709 25002
rect 15775 24970 15809 25002
rect 15875 24970 15909 25002
rect 15375 24870 15409 24904
rect 15475 24870 15509 24904
rect 15575 24870 15609 24904
rect 15675 24870 15709 24904
rect 15775 24870 15809 24904
rect 15875 24870 15909 24904
rect 15375 24770 15409 24804
rect 15475 24770 15509 24804
rect 15575 24770 15609 24804
rect 15675 24770 15709 24804
rect 15775 24770 15809 24804
rect 15875 24770 15909 24804
rect 15375 24676 15409 24704
rect 15375 24670 15381 24676
rect 15381 24670 15409 24676
rect 15475 24670 15509 24704
rect 15575 24670 15609 24704
rect 15675 24676 15709 24704
rect 15775 24676 15809 24704
rect 15875 24676 15909 24704
rect 15675 24670 15707 24676
rect 15707 24670 15709 24676
rect 15775 24670 15797 24676
rect 15797 24670 15809 24676
rect 15875 24670 15887 24676
rect 15887 24670 15909 24676
rect 16092 25245 16097 25279
rect 16097 25278 16508 25279
rect 16097 25245 16211 25278
rect 16092 25244 16211 25245
rect 16211 25244 16245 25278
rect 16245 25244 16368 25278
rect 16368 25244 16402 25278
rect 16402 25244 16508 25278
rect 17424 25334 17555 25368
rect 17555 25334 17589 25368
rect 17589 25334 17590 25368
rect 17424 25279 17590 25334
rect 16092 25189 16508 25244
rect 16092 25155 16097 25189
rect 16097 25188 16508 25189
rect 16097 25155 16211 25188
rect 16092 25154 16211 25155
rect 16211 25154 16245 25188
rect 16245 25154 16368 25188
rect 16368 25154 16402 25188
rect 16402 25154 16508 25188
rect 16092 25105 16508 25154
rect 16088 24705 16097 24712
rect 16097 24705 16211 24712
rect 16088 24704 16211 24705
rect 16211 24704 16245 24712
rect 16245 24704 16368 24712
rect 16368 24704 16402 24712
rect 16402 24704 16530 24712
rect 16088 24668 16530 24704
rect 16088 24649 16517 24668
rect 16088 24615 16097 24649
rect 16097 24648 16517 24649
rect 16097 24615 16211 24648
rect 14743 24559 15173 24578
rect 14743 24525 14753 24559
rect 14753 24558 15173 24559
rect 14753 24525 14867 24558
rect 14743 24524 14867 24525
rect 14867 24524 14901 24558
rect 14901 24524 15024 24558
rect 15024 24524 15058 24558
rect 15058 24544 15173 24558
rect 15173 24544 15185 24578
rect 15058 24524 15185 24544
rect 14743 24496 15185 24524
rect 16088 24614 16211 24615
rect 16211 24614 16245 24648
rect 16245 24614 16368 24648
rect 16368 24614 16402 24648
rect 16402 24634 16517 24648
rect 16517 24634 16530 24668
rect 16402 24614 16530 24634
rect 16088 24578 16530 24614
rect 16719 25182 16725 25204
rect 16725 25182 16753 25204
rect 16719 25170 16753 25182
rect 16819 25170 16853 25204
rect 16919 25170 16953 25204
rect 17019 25182 17051 25204
rect 17051 25182 17053 25204
rect 17119 25182 17141 25204
rect 17141 25182 17153 25204
rect 17219 25182 17231 25204
rect 17231 25182 17253 25204
rect 17019 25170 17053 25182
rect 17119 25170 17153 25182
rect 17219 25170 17253 25182
rect 16719 25092 16725 25104
rect 16725 25092 16753 25104
rect 16719 25070 16753 25092
rect 16819 25070 16853 25104
rect 16919 25070 16953 25104
rect 17019 25092 17051 25104
rect 17051 25092 17053 25104
rect 17119 25092 17141 25104
rect 17141 25092 17153 25104
rect 17219 25092 17231 25104
rect 17231 25092 17253 25104
rect 17019 25070 17053 25092
rect 17119 25070 17153 25092
rect 17219 25070 17253 25092
rect 16719 25002 16725 25004
rect 16725 25002 16753 25004
rect 16719 24970 16753 25002
rect 16819 24970 16853 25004
rect 16919 24970 16953 25004
rect 17019 25002 17051 25004
rect 17051 25002 17053 25004
rect 17119 25002 17141 25004
rect 17141 25002 17153 25004
rect 17219 25002 17231 25004
rect 17231 25002 17253 25004
rect 17019 24970 17053 25002
rect 17119 24970 17153 25002
rect 17219 24970 17253 25002
rect 16719 24870 16753 24904
rect 16819 24870 16853 24904
rect 16919 24870 16953 24904
rect 17019 24870 17053 24904
rect 17119 24870 17153 24904
rect 17219 24870 17253 24904
rect 16719 24770 16753 24804
rect 16819 24770 16853 24804
rect 16919 24770 16953 24804
rect 17019 24770 17053 24804
rect 17119 24770 17153 24804
rect 17219 24770 17253 24804
rect 16719 24676 16753 24704
rect 16719 24670 16725 24676
rect 16725 24670 16753 24676
rect 16819 24670 16853 24704
rect 16919 24670 16953 24704
rect 17019 24676 17053 24704
rect 17119 24676 17153 24704
rect 17219 24676 17253 24704
rect 17019 24670 17051 24676
rect 17051 24670 17053 24676
rect 17119 24670 17141 24676
rect 17141 24670 17153 24676
rect 17219 24670 17231 24676
rect 17231 24670 17253 24676
rect 17424 25245 17441 25279
rect 17441 25278 17590 25279
rect 17441 25245 17555 25278
rect 17424 25244 17555 25245
rect 17555 25244 17589 25278
rect 17589 25244 17590 25278
rect 17424 25189 17590 25244
rect 17424 25155 17441 25189
rect 17441 25188 17590 25189
rect 17441 25155 17555 25188
rect 17424 25154 17555 25155
rect 17555 25154 17589 25188
rect 17589 25154 17590 25188
rect 17424 25099 17590 25154
rect 17424 25065 17441 25099
rect 17441 25098 17590 25099
rect 17441 25065 17555 25098
rect 17424 25064 17555 25065
rect 17555 25064 17589 25098
rect 17589 25064 17590 25098
rect 17424 25009 17590 25064
rect 17424 24975 17441 25009
rect 17441 25008 17590 25009
rect 17441 24975 17555 25008
rect 17424 24974 17555 24975
rect 17555 24974 17589 25008
rect 17589 24974 17590 25008
rect 17424 24919 17590 24974
rect 17424 24885 17441 24919
rect 17441 24918 17590 24919
rect 17441 24885 17555 24918
rect 17424 24884 17555 24885
rect 17555 24884 17589 24918
rect 17589 24884 17590 24918
rect 17424 24829 17590 24884
rect 17424 24795 17441 24829
rect 17441 24828 17590 24829
rect 17441 24795 17555 24828
rect 17424 24794 17555 24795
rect 17555 24794 17589 24828
rect 17589 24794 17590 24828
rect 17424 24739 17590 24794
rect 17424 24705 17441 24739
rect 17441 24738 17590 24739
rect 17441 24705 17555 24738
rect 17424 24704 17555 24705
rect 17555 24704 17589 24738
rect 17589 24704 17590 24738
rect 17424 24649 17590 24704
rect 17424 24615 17441 24649
rect 17441 24648 17590 24649
rect 17441 24615 17555 24648
rect 16088 24559 16517 24578
rect 16088 24525 16097 24559
rect 16097 24558 16517 24559
rect 16097 24525 16211 24558
rect 16088 24524 16211 24525
rect 16211 24524 16245 24558
rect 16245 24524 16368 24558
rect 16368 24524 16402 24558
rect 16402 24544 16517 24558
rect 16517 24544 16530 24578
rect 16402 24524 16530 24544
rect 16088 24496 16530 24524
rect 17424 24614 17555 24615
rect 17555 24614 17589 24648
rect 17589 24614 17590 24648
rect 17424 24559 17590 24614
rect 17424 24525 17441 24559
rect 17441 24558 17590 24559
rect 17441 24525 17555 24558
rect 17424 24524 17555 24525
rect 17555 24524 17589 24558
rect 17589 24524 17590 24558
rect 17424 24496 17590 24524
rect 5742 24468 13887 24496
rect 13887 24468 13921 24496
rect 13921 24468 13977 24496
rect 13977 24468 14011 24496
rect 14011 24468 14067 24496
rect 14067 24468 14101 24496
rect 14101 24468 14157 24496
rect 14157 24468 14191 24496
rect 14191 24468 14247 24496
rect 14247 24468 14281 24496
rect 14281 24468 14337 24496
rect 14337 24468 14371 24496
rect 14371 24468 14427 24496
rect 14427 24468 14461 24496
rect 14461 24468 14517 24496
rect 14517 24468 14551 24496
rect 14551 24468 14607 24496
rect 14607 24468 14641 24496
rect 14641 24468 15231 24496
rect 15231 24468 15265 24496
rect 15265 24468 15321 24496
rect 15321 24468 15355 24496
rect 15355 24468 15411 24496
rect 15411 24468 15445 24496
rect 15445 24468 15501 24496
rect 15501 24468 15535 24496
rect 15535 24468 15591 24496
rect 15591 24468 15625 24496
rect 15625 24468 15681 24496
rect 15681 24468 15715 24496
rect 15715 24468 15771 24496
rect 15771 24468 15805 24496
rect 15805 24468 15861 24496
rect 15861 24468 15895 24496
rect 15895 24468 15951 24496
rect 15951 24468 15985 24496
rect 15985 24468 16575 24496
rect 16575 24468 16609 24496
rect 16609 24468 16665 24496
rect 16665 24468 16699 24496
rect 16699 24468 16755 24496
rect 16755 24468 16789 24496
rect 16789 24468 16845 24496
rect 16845 24468 16879 24496
rect 16879 24468 16935 24496
rect 16935 24468 16969 24496
rect 16969 24468 17025 24496
rect 17025 24468 17059 24496
rect 17059 24468 17115 24496
rect 17115 24468 17149 24496
rect 17149 24468 17205 24496
rect 17205 24468 17239 24496
rect 17239 24468 17295 24496
rect 17295 24468 17329 24496
rect 17329 24468 17592 24496
rect 5742 24434 13680 24468
rect 13680 24434 13714 24468
rect 13714 24434 14867 24468
rect 14867 24434 14901 24468
rect 14901 24434 15024 24468
rect 15024 24434 15058 24468
rect 15058 24434 16211 24468
rect 16211 24434 16245 24468
rect 16245 24434 16368 24468
rect 16368 24434 16402 24468
rect 16402 24434 17555 24468
rect 17555 24434 17589 24468
rect 17589 24434 17592 24468
rect 5742 24387 17592 24434
rect 5742 24378 17598 24387
rect 5742 24344 13680 24378
rect 13680 24344 13714 24378
rect 13714 24355 14867 24378
rect 13714 24344 13781 24355
rect 5742 24321 13781 24344
rect 13781 24321 13815 24355
rect 13815 24321 13871 24355
rect 13871 24321 13905 24355
rect 13905 24321 13961 24355
rect 13961 24321 13995 24355
rect 13995 24321 14051 24355
rect 14051 24321 14085 24355
rect 14085 24321 14141 24355
rect 14141 24321 14175 24355
rect 14175 24321 14231 24355
rect 14231 24321 14265 24355
rect 14265 24321 14321 24355
rect 14321 24321 14355 24355
rect 14355 24321 14411 24355
rect 14411 24321 14445 24355
rect 14445 24321 14501 24355
rect 14501 24321 14535 24355
rect 14535 24321 14591 24355
rect 14591 24321 14625 24355
rect 14625 24321 14681 24355
rect 14681 24321 14715 24355
rect 14715 24321 14771 24355
rect 14771 24321 14805 24355
rect 14805 24344 14867 24355
rect 14867 24344 14901 24378
rect 14901 24344 15024 24378
rect 15024 24344 15058 24378
rect 15058 24355 16211 24378
rect 15058 24344 15125 24355
rect 14805 24321 15125 24344
rect 15125 24321 15159 24355
rect 15159 24321 15215 24355
rect 15215 24321 15249 24355
rect 15249 24321 15305 24355
rect 15305 24321 15339 24355
rect 15339 24321 15395 24355
rect 15395 24321 15429 24355
rect 15429 24321 15485 24355
rect 15485 24321 15519 24355
rect 15519 24321 15575 24355
rect 15575 24321 15609 24355
rect 15609 24321 15665 24355
rect 15665 24321 15699 24355
rect 15699 24321 15755 24355
rect 15755 24321 15789 24355
rect 15789 24321 15845 24355
rect 15845 24321 15879 24355
rect 15879 24321 15935 24355
rect 15935 24321 15969 24355
rect 15969 24321 16025 24355
rect 16025 24321 16059 24355
rect 16059 24321 16115 24355
rect 16115 24321 16149 24355
rect 16149 24344 16211 24355
rect 16211 24344 16245 24378
rect 16245 24344 16368 24378
rect 16368 24344 16402 24378
rect 16402 24355 17555 24378
rect 16402 24344 16469 24355
rect 16149 24321 16469 24344
rect 16469 24321 16503 24355
rect 16503 24321 16559 24355
rect 16559 24321 16593 24355
rect 16593 24321 16649 24355
rect 16649 24321 16683 24355
rect 16683 24321 16739 24355
rect 16739 24321 16773 24355
rect 16773 24321 16829 24355
rect 16829 24321 16863 24355
rect 16863 24321 16919 24355
rect 16919 24321 16953 24355
rect 16953 24321 17009 24355
rect 17009 24321 17043 24355
rect 17043 24321 17099 24355
rect 17099 24321 17133 24355
rect 17133 24321 17189 24355
rect 17189 24321 17223 24355
rect 17223 24321 17279 24355
rect 17279 24321 17313 24355
rect 17313 24321 17369 24355
rect 17369 24321 17403 24355
rect 17403 24321 17459 24355
rect 17459 24321 17493 24355
rect 17493 24344 17555 24355
rect 17555 24344 17589 24378
rect 17589 24344 17598 24378
rect 17493 24321 17598 24344
rect 5742 24236 17598 24321
rect 5742 24202 6038 24236
rect 6038 24202 6366 24236
rect 6366 24202 6524 24236
rect 6524 24202 6852 24236
rect 6852 24202 7010 24236
rect 7010 24202 7338 24236
rect 7338 24202 7496 24236
rect 7496 24202 7824 24236
rect 7824 24202 7982 24236
rect 7982 24202 8310 24236
rect 8310 24202 8468 24236
rect 8468 24202 8796 24236
rect 8796 24202 8954 24236
rect 8954 24202 9282 24236
rect 9282 24202 9440 24236
rect 9440 24202 9768 24236
rect 9768 24202 9926 24236
rect 9926 24202 10254 24236
rect 10254 24202 10412 24236
rect 10412 24202 10740 24236
rect 10740 24211 17598 24236
rect 10740 24202 11232 24211
rect 13517 24204 17598 24211
rect 5742 24198 11232 24202
rect 5742 24140 5981 24198
rect 5742 19972 5942 24140
rect 5942 19972 5976 24140
rect 5976 19972 5981 24140
rect 6428 24140 6462 24198
rect 6164 24068 6240 24102
rect 6080 20072 6114 24040
rect 6290 20072 6324 24040
rect 6164 20010 6240 20044
rect 5742 19954 5981 19972
rect 6428 19972 6462 24140
rect 6914 24140 6948 24198
rect 6650 24068 6726 24102
rect 6566 20072 6600 24040
rect 6776 20072 6810 24040
rect 6650 20010 6726 20044
rect 6428 19954 6462 19972
rect 6914 19972 6948 24140
rect 7400 24140 7434 24198
rect 7136 24068 7212 24102
rect 7052 20072 7086 24040
rect 7262 20072 7296 24040
rect 7136 20010 7212 20044
rect 6914 19954 6948 19972
rect 7400 19972 7434 24140
rect 7886 24140 7920 24198
rect 7622 24068 7698 24102
rect 7538 20072 7572 24040
rect 7748 20072 7782 24040
rect 7622 20010 7698 20044
rect 7400 19954 7434 19972
rect 7886 19972 7920 24140
rect 8372 24140 8406 24198
rect 8108 24068 8184 24102
rect 8024 20072 8058 24040
rect 8234 20072 8268 24040
rect 8108 20010 8184 20044
rect 7886 19954 7920 19972
rect 8372 19972 8406 24140
rect 8858 24140 8892 24198
rect 8594 24068 8670 24102
rect 8510 20072 8544 24040
rect 8720 20072 8754 24040
rect 8594 20010 8670 20044
rect 8372 19954 8406 19972
rect 8858 19972 8892 24140
rect 9344 24140 9378 24198
rect 9080 24068 9156 24102
rect 8996 20072 9030 24040
rect 9206 20072 9240 24040
rect 9080 20010 9156 20044
rect 8858 19954 8892 19972
rect 9344 19972 9378 24140
rect 9830 24140 9864 24198
rect 9566 24068 9642 24102
rect 9482 20072 9516 24040
rect 9692 20072 9726 24040
rect 9566 20010 9642 20044
rect 9344 19954 9378 19972
rect 9830 19972 9864 24140
rect 10316 24140 10350 24198
rect 10052 24068 10128 24102
rect 9968 20072 10002 24040
rect 10178 20072 10212 24040
rect 10052 20010 10128 20044
rect 9830 19954 9864 19972
rect 10316 19972 10350 24140
rect 10538 24068 10614 24102
rect 10454 20072 10488 24040
rect 10664 20072 10698 24040
rect 10538 20010 10614 20044
rect 10316 19954 10350 19972
rect 10771 24140 10855 24198
rect 10771 19972 10802 24140
rect 10802 19972 10836 24140
rect 10836 23510 10855 24140
rect 15561 24049 17598 24204
rect 15561 23843 20149 24049
rect 15564 23829 20149 23843
rect 15564 23795 15759 23829
rect 15759 23795 19927 23829
rect 19927 23795 20149 23829
rect 15564 23789 20149 23795
rect 10836 23429 15595 23510
rect 10836 23395 11303 23429
rect 11303 23395 15471 23429
rect 15471 23395 15595 23429
rect 10836 23364 15595 23395
rect 10836 23363 10918 23364
rect 10836 20784 10855 23363
rect 11074 23333 11220 23364
rect 11074 22505 11207 23333
rect 11207 22505 11220 23333
rect 11403 23257 15371 23291
rect 11341 22631 11375 23207
rect 15399 22631 15433 23207
rect 11403 22547 15371 22581
rect 11074 22356 11220 22505
rect 19965 23733 20149 23789
rect 15859 23657 19827 23691
rect 15797 22631 15831 23607
rect 19855 22631 19889 23607
rect 15859 22547 19827 22581
rect 19965 22505 19989 23733
rect 19989 22505 20023 23733
rect 20023 22505 20149 23733
rect 19965 22387 20149 22505
rect 11074 22337 15126 22356
rect 11080 22172 15126 22337
rect 11200 22061 11261 22172
rect 16147 22157 20149 22387
rect 16147 22146 19927 22157
rect 19927 22146 20149 22157
rect 11200 20833 11214 22061
rect 11214 20833 11248 22061
rect 11248 20833 11261 22061
rect 11410 21985 15378 22019
rect 11348 20959 11382 21935
rect 15406 20959 15440 21935
rect 15530 21161 15540 21768
rect 11410 20875 15378 20909
rect 11200 20784 11261 20833
rect 15532 20833 15540 21161
rect 15540 20833 15574 21768
rect 15574 21233 15663 21768
rect 15663 21233 15686 21768
rect 19965 22061 20149 22146
rect 15859 21985 19827 22019
rect 15797 21359 15831 21935
rect 19855 21359 19889 21935
rect 15859 21275 19827 21309
rect 15574 21189 15686 21233
rect 19965 21233 19989 22061
rect 19989 21233 20023 22061
rect 20023 21233 20149 22061
rect 19965 21189 20149 21233
rect 15574 21171 20149 21189
rect 15574 21137 15759 21171
rect 15759 21137 19927 21171
rect 19927 21137 20149 21171
rect 15574 21081 20149 21137
rect 15574 20833 15600 21081
rect 10836 20783 11263 20784
rect 15532 20783 15600 20833
rect 10836 20771 15603 20783
rect 10836 20737 11310 20771
rect 11310 20737 15478 20771
rect 15478 20737 15603 20771
rect 10836 20696 15603 20737
rect 10836 19972 10855 20696
rect 10771 19954 10855 19972
rect 5742 19910 10855 19954
rect 5742 19876 6038 19910
rect 6038 19876 6366 19910
rect 6366 19876 6524 19910
rect 6524 19876 6852 19910
rect 6852 19876 7010 19910
rect 7010 19876 7338 19910
rect 7338 19876 7496 19910
rect 7496 19876 7824 19910
rect 7824 19876 7982 19910
rect 7982 19876 8310 19910
rect 8310 19876 8468 19910
rect 8468 19876 8796 19910
rect 8796 19876 8954 19910
rect 8954 19876 9282 19910
rect 9282 19876 9440 19910
rect 9440 19876 9768 19910
rect 9768 19876 9926 19910
rect 9926 19876 10254 19910
rect 10254 19876 10412 19910
rect 10412 19876 10740 19910
rect 10740 19876 10855 19910
rect 5742 19739 10855 19876
rect 5742 19731 10825 19739
rect 6141 19270 20095 19366
rect 6141 19246 6320 19270
rect 6320 19246 10488 19270
rect 10488 19246 11408 19270
rect 11408 19246 15576 19270
rect 15576 19246 15734 19270
rect 15734 19246 19902 19270
rect 19902 19246 20095 19270
rect 6141 19174 6252 19246
rect 6141 18092 6224 19174
rect 6224 18092 6252 19174
rect 10574 19174 11339 19246
rect 6420 19098 10388 19132
rect 6358 18763 6392 19039
rect 10416 18763 10450 19039
rect 6420 18670 10388 18704
rect 6420 18562 10388 18596
rect 6358 18227 6392 18503
rect 10416 18227 10450 18503
rect 6420 18134 10388 18168
rect 6141 17774 6252 18092
rect 10574 18092 10584 19174
rect 10584 18092 11312 19174
rect 6141 16928 6224 17774
rect 6224 16928 6252 17774
rect 10574 17774 11312 18092
rect 6420 17698 10388 17732
rect 6358 17063 6392 17639
rect 10416 17063 10450 17639
rect 6420 16970 10388 17004
rect 6141 16875 6252 16928
rect 10574 16928 10584 17774
rect 10584 16928 11312 17774
rect 11312 16928 11339 19174
rect 11508 19098 15476 19132
rect 11446 17063 11480 19039
rect 15504 17063 15538 19039
rect 11508 16970 15476 17004
rect 10574 16875 11339 16928
rect 6136 16866 11339 16875
rect 19971 19174 20095 19246
rect 15834 19098 19802 19132
rect 15772 17063 15806 19039
rect 19830 17063 19864 19039
rect 15834 16970 19802 17004
rect 19971 18903 19998 19174
rect 19998 18983 20095 19174
rect 20576 18983 21831 18992
rect 19989 16928 19998 18903
rect 19998 18902 21831 18983
rect 19998 18868 20776 18902
rect 20776 18868 21122 18902
rect 21122 18868 21280 18902
rect 21280 18868 21626 18902
rect 21626 18868 21831 18902
rect 19998 18859 21831 18868
rect 19998 18806 20718 18859
rect 19998 16928 20680 18806
rect 6136 16832 6320 16866
rect 6320 16832 10488 16866
rect 10488 16832 11339 16866
rect 6136 16770 11339 16832
rect 6136 16741 11312 16770
rect 8056 15066 11312 16741
rect 8056 15041 8330 15066
rect 8330 15041 10488 15066
rect 10488 15041 11312 15066
rect 8056 14970 8243 15041
rect 8056 14524 8234 14970
rect 8234 14524 8243 14970
rect 10574 14970 11312 15041
rect 8430 14894 10388 14928
rect 8368 14659 8402 14835
rect 10416 14659 10450 14835
rect 8430 14566 10388 14600
rect 8056 14464 8243 14524
rect 10574 14524 10584 14970
rect 10584 14524 11312 14970
rect 11312 14524 11339 16770
rect 11508 16694 15476 16728
rect 11446 14659 11480 16635
rect 15504 14659 15538 16635
rect 11508 14566 15476 14600
rect 10574 14464 11339 14524
rect 19989 16770 20680 16928
rect 15834 16694 19802 16728
rect 15772 14659 15806 16635
rect 19830 14659 19864 16635
rect 15834 14566 19802 14600
rect 19989 14524 19998 16770
rect 19998 14638 20680 16770
rect 20680 14638 20714 18806
rect 20714 14638 20718 18806
rect 19998 14524 20718 14638
rect 20911 18734 20987 18768
rect 20818 14738 20852 18706
rect 21046 14738 21080 18706
rect 20911 14676 20987 14710
rect 21415 18734 21491 18768
rect 21322 14738 21356 18706
rect 21550 14738 21584 18706
rect 21415 14676 21491 14710
rect 21688 18806 21822 18859
rect 21688 14638 21722 18806
rect 21722 14638 21822 18806
rect 19989 14464 20718 14524
rect 21688 14464 21822 14638
rect 8056 14462 21822 14464
rect 8056 14428 8330 14462
rect 8330 14428 10488 14462
rect 10488 14428 11408 14462
rect 11408 14428 15576 14462
rect 15576 14428 15734 14462
rect 15734 14428 19902 14462
rect 19902 14428 21822 14462
rect 8056 14418 21822 14428
rect 8056 14001 21806 14418
rect 7800 12663 10778 12824
rect 7800 12572 10779 12663
rect 7796 12542 10779 12572
rect 7796 12519 8035 12542
rect 8035 12519 10213 12542
rect 10213 12519 10779 12542
rect 7796 12446 7999 12519
rect 7796 12000 7939 12446
rect 7939 12000 7973 12446
rect 7973 12000 7999 12446
rect 7796 11969 7999 12000
rect 10284 12446 10779 12519
rect 8135 12370 10113 12404
rect 8073 12135 8107 12311
rect 10141 12135 10175 12311
rect 8135 12042 10113 12076
rect 10284 12000 10309 12446
rect 10309 12000 10779 12446
rect 10284 11969 10779 12000
rect 5840 11938 10779 11969
rect 5840 11904 8035 11938
rect 8035 11904 10213 11938
rect 10213 11904 10779 11938
rect 5840 11779 10779 11904
rect 5840 11757 6035 11779
rect 6035 11757 10203 11779
rect 10203 11757 10779 11779
rect 5840 11683 5983 11757
rect 5840 11037 5939 11683
rect 5939 11037 5973 11683
rect 5973 11037 5983 11683
rect 5840 10982 5983 11037
rect 10284 11683 10779 11757
rect 6135 11607 10103 11641
rect 6073 11172 6107 11548
rect 10131 11172 10165 11548
rect 6135 11079 10103 11113
rect 10284 11037 10299 11683
rect 10299 11037 10779 11683
rect 10284 10982 10779 11037
rect 5840 10975 10779 10982
rect 5840 10941 6035 10975
rect 6035 10941 10203 10975
rect 10203 10941 10779 10975
rect 5840 10811 10779 10941
rect 5840 10801 9013 10811
rect 9013 10801 9661 10811
rect 9661 10801 9945 10811
rect 9945 10806 10593 10811
rect 10593 10806 10779 10811
rect 9945 10801 10361 10806
rect 5844 10697 6065 10801
rect 5844 9951 6051 10697
rect 6051 9951 6065 10697
rect 6247 10621 6695 10655
rect 6185 10086 6219 10562
rect 6723 10086 6757 10562
rect 6247 9993 6695 10027
rect 5844 9655 6065 9951
rect 7183 10621 7631 10655
rect 7121 10086 7155 10562
rect 7659 10086 7693 10562
rect 7183 9993 7631 10027
rect 7787 10697 7942 10801
rect 7787 9951 7793 10697
rect 7793 9951 7827 10697
rect 7827 9951 7942 10697
rect 5844 8909 6051 9655
rect 6051 8909 6065 9655
rect 6247 9579 6695 9613
rect 6185 9044 6219 9520
rect 6723 9044 6757 9520
rect 6247 8951 6695 8985
rect 5844 8871 6065 8909
rect 7183 9579 7631 9613
rect 7121 9044 7155 9520
rect 7659 9044 7693 9520
rect 7183 8951 7631 8985
rect 7787 9655 7942 9951
rect 7787 8909 7793 9655
rect 7793 8909 7827 9655
rect 7827 8909 7942 9655
rect 7787 8871 7942 8909
rect 8812 10715 8950 10801
rect 8812 9969 8917 10715
rect 8917 9969 8950 10715
rect 9113 10639 9561 10673
rect 9051 10104 9085 10580
rect 9589 10104 9623 10580
rect 9113 10011 9561 10045
rect 8812 9630 8950 9969
rect 10045 10639 10493 10673
rect 9983 10104 10017 10580
rect 10521 10104 10555 10580
rect 10045 10011 10493 10045
rect 10655 10715 10776 10806
rect 10655 9969 10689 10715
rect 10689 9969 10776 10715
rect 8812 8884 8917 9630
rect 8917 8884 8950 9630
rect 9113 9554 9561 9588
rect 9051 9019 9085 9495
rect 9589 9019 9623 9495
rect 9113 8926 9561 8960
rect 10045 9554 10493 9588
rect 9983 9019 10017 9495
rect 10521 9019 10555 9495
rect 10045 8926 10493 8960
rect 5844 8847 7960 8871
rect 5844 8813 6147 8847
rect 6147 8813 6795 8847
rect 6795 8813 7083 8847
rect 7083 8813 7731 8847
rect 7731 8813 7960 8847
rect 5844 8767 7960 8813
rect 8812 8863 8950 8884
rect 10655 9630 10776 9969
rect 10655 8884 10689 9630
rect 10689 8884 10776 9630
rect 10655 8863 10776 8884
rect 8812 8822 10776 8863
rect 8812 8788 9013 8822
rect 9013 8788 9661 8822
rect 9661 8788 9945 8822
rect 9945 8788 10593 8822
rect 10593 8788 10776 8822
rect 8812 8741 10776 8788
rect 11880 11114 12899 11117
rect 11848 11079 12899 11114
rect 11848 11049 12901 11079
rect 11848 11015 11973 11049
rect 11973 11015 12757 11049
rect 12757 11015 12901 11049
rect 11848 11006 12901 11015
rect 11848 10989 11967 11006
rect 11848 10533 11913 10989
rect 11913 10533 11947 10989
rect 11947 10533 11967 10989
rect 11848 10404 11967 10533
rect 12095 10912 12163 10946
rect 12253 10912 12321 10946
rect 12411 10912 12479 10946
rect 12569 10912 12637 10946
rect 12033 10677 12067 10853
rect 12191 10677 12225 10853
rect 12349 10677 12383 10853
rect 12507 10677 12541 10853
rect 12665 10677 12699 10853
rect 12095 10584 12163 10618
rect 12253 10584 12321 10618
rect 12411 10584 12479 10618
rect 12569 10584 12637 10618
rect 12773 10989 12901 11006
rect 12773 10533 12783 10989
rect 12783 10533 12817 10989
rect 12817 10533 12901 10989
rect 12773 10418 12901 10533
rect 13753 10853 20417 11042
rect 11241 9764 11310 9898
rect 11241 9336 11283 9764
rect 11283 9336 11310 9764
rect 11723 9764 11848 9898
rect 11479 9688 11547 9722
rect 11417 9462 11451 9638
rect 11575 9462 11609 9638
rect 11479 9378 11547 9412
rect 11241 9287 11310 9336
rect 11723 9336 11743 9764
rect 11743 9336 11839 9764
rect 11839 9336 11848 9764
rect 12280 9764 12405 9901
rect 12035 9688 12103 9722
rect 11973 9462 12007 9638
rect 12131 9462 12165 9638
rect 12035 9378 12103 9412
rect 11723 9287 11848 9336
rect 12280 9336 12299 9764
rect 12299 9336 12395 9764
rect 12395 9336 12405 9764
rect 12844 9764 12969 9893
rect 12591 9688 12659 9722
rect 12529 9462 12563 9638
rect 12687 9462 12721 9638
rect 12591 9378 12659 9412
rect 12280 9287 12405 9336
rect 12844 9336 12855 9764
rect 12855 9336 12951 9764
rect 12951 9336 12969 9764
rect 13384 9764 13448 9900
rect 13147 9688 13215 9722
rect 13085 9462 13119 9638
rect 13243 9462 13277 9638
rect 13147 9378 13215 9412
rect 12844 9287 12969 9336
rect 13384 9336 13411 9764
rect 13411 9336 13448 9764
rect 13384 9287 13448 9336
rect 11241 9274 13446 9287
rect 11241 9240 11379 9274
rect 11379 9240 11647 9274
rect 11647 9240 11935 9274
rect 11935 9240 12203 9274
rect 12203 9240 12491 9274
rect 12491 9240 12759 9274
rect 12759 9240 13047 9274
rect 13047 9240 13315 9274
rect 13315 9240 13446 9274
rect 11241 9173 13446 9240
rect 8821 8737 10776 8741
rect 10655 8728 10776 8737
rect 8523 8640 8589 8650
rect 5318 8630 8589 8640
rect 5295 8626 8589 8630
rect 5295 8610 10790 8626
rect 5295 8609 9985 8610
rect 5295 8575 5427 8609
rect 5427 8575 6795 8609
rect 6795 8575 7083 8609
rect 7083 8575 8451 8609
rect 8451 8575 9013 8609
rect 9013 8575 9621 8609
rect 9621 8576 9985 8609
rect 9985 8576 10593 8610
rect 10593 8576 10790 8610
rect 9621 8575 10790 8576
rect 5295 8564 10790 8575
rect 5295 8560 8589 8564
rect 5295 8513 5375 8560
rect 5295 8085 5331 8513
rect 5331 8085 5365 8513
rect 5365 8085 5375 8513
rect 5295 8009 5375 8085
rect 5527 8437 6695 8471
rect 5465 8211 5499 8387
rect 6723 8211 6757 8387
rect 5527 8127 6695 8161
rect 8523 8513 8589 8560
rect 7183 8437 8351 8471
rect 7121 8211 7155 8387
rect 8379 8211 8413 8387
rect 7183 8127 8351 8161
rect 8523 8085 8547 8513
rect 8547 8085 8589 8513
rect 8523 8009 8589 8085
rect 5295 7989 5427 8009
rect 5427 7989 6795 8009
rect 6795 7989 7083 8009
rect 7083 7989 8451 8009
rect 8451 7995 8589 8009
rect 8824 8513 8961 8564
rect 8824 8085 8917 8513
rect 8917 8085 8951 8513
rect 8951 8085 8961 8513
rect 8824 7995 8961 8085
rect 9704 8514 9897 8564
rect 9704 8513 9889 8514
rect 9113 8437 9521 8471
rect 9051 8211 9085 8387
rect 9549 8211 9583 8387
rect 9113 8127 9521 8161
rect 9704 8085 9717 8513
rect 9717 8086 9889 8513
rect 9889 8086 9897 8514
rect 10665 8514 10790 8564
rect 10085 8438 10493 8472
rect 10023 8212 10057 8388
rect 10521 8212 10555 8388
rect 10085 8128 10493 8162
rect 9717 8085 9897 8086
rect 9704 7995 9897 8085
rect 10665 8086 10689 8514
rect 10689 8086 10790 8514
rect 10665 7995 10790 8086
rect 8451 7989 9013 7995
rect 9013 7989 9621 7995
rect 9621 7990 9985 7995
rect 9985 7990 10593 7995
rect 10593 7990 10802 7995
rect 9621 7989 10802 7990
rect 5295 7933 10802 7989
rect 5295 7893 8589 7933
rect 5295 7869 5427 7893
rect 5427 7869 6795 7893
rect 6795 7869 7083 7893
rect 7083 7869 8451 7893
rect 8451 7869 8589 7893
rect 5295 7797 5375 7869
rect 5295 7369 5331 7797
rect 5331 7369 5365 7797
rect 5365 7369 5375 7797
rect 5295 7295 5375 7369
rect 5527 7721 6695 7755
rect 5465 7495 5499 7671
rect 6723 7495 6757 7671
rect 5527 7411 6695 7445
rect 8523 7797 8589 7869
rect 7183 7721 8351 7755
rect 7121 7495 7155 7671
rect 8379 7495 8413 7671
rect 7183 7411 8351 7445
rect 8523 7369 8547 7797
rect 8547 7369 8589 7797
rect 8523 7295 8589 7369
rect 5295 7273 5427 7295
rect 5427 7273 6795 7295
rect 6795 7273 7083 7295
rect 7083 7273 8451 7295
rect 8451 7273 8589 7295
rect 5295 7177 8589 7273
rect 5295 7155 5427 7177
rect 5427 7155 6795 7177
rect 6795 7155 7083 7177
rect 7083 7155 8451 7177
rect 8451 7155 8589 7177
rect 5295 7081 5375 7155
rect 5295 6653 5331 7081
rect 5331 6653 5365 7081
rect 5365 6653 5375 7081
rect 5295 6564 5375 6653
rect 5527 7005 6695 7039
rect 5465 6779 5499 6955
rect 6723 6779 6757 6955
rect 5527 6695 6695 6729
rect 8523 7081 8589 7155
rect 7183 7005 8351 7039
rect 7121 6779 7155 6955
rect 8379 6779 8413 6955
rect 7183 6695 8351 6729
rect 8523 6653 8547 7081
rect 8547 6653 8589 7081
rect 8523 6564 8589 6653
rect 5295 6557 5427 6564
rect 5427 6557 6795 6564
rect 6795 6557 7083 6564
rect 7083 6557 8451 6564
rect 8451 6557 8589 6564
rect 5295 6461 8589 6557
rect 5295 6427 5427 6461
rect 5427 6427 6795 6461
rect 6795 6427 7083 6461
rect 7083 6427 8451 6461
rect 8451 6427 8589 6461
rect 5295 6424 8589 6427
rect 5295 6365 5375 6424
rect 5295 5937 5331 6365
rect 5331 5937 5365 6365
rect 5365 5937 5375 6365
rect 5295 5867 5375 5937
rect 5527 6289 6695 6323
rect 5465 6063 5499 6239
rect 6723 6063 6757 6239
rect 5527 5979 6695 6013
rect 8523 6365 8589 6424
rect 7183 6289 8351 6323
rect 7121 6063 7155 6239
rect 8379 6063 8413 6239
rect 7183 5979 8351 6013
rect 8523 5937 8547 6365
rect 8547 5937 8589 6365
rect 8523 5867 8589 5937
rect 5295 5841 5427 5867
rect 5427 5841 6795 5867
rect 6795 5841 7083 5867
rect 7083 5841 8451 5867
rect 8451 5841 8589 5867
rect 5295 5730 8589 5841
rect 5335 5727 8589 5730
rect 8523 5720 8589 5727
rect 13753 2391 13873 10853
rect 14113 10282 14151 10679
rect 14113 6783 14151 7180
rect 14409 10282 14447 10679
rect 14409 6783 14447 7180
rect 14705 10282 14743 10679
rect 14705 6783 14743 7180
rect 15001 10282 15039 10679
rect 15001 6783 15039 7180
rect 15297 10282 15335 10679
rect 15297 6783 15335 7180
rect 15593 10282 15631 10679
rect 15593 6783 15631 7180
rect 15889 10282 15927 10679
rect 15889 6783 15927 7180
rect 16185 10282 16223 10679
rect 16185 6783 16223 7180
rect 16585 10277 20388 10288
rect 16585 10100 20400 10277
rect 16671 9726 16739 9760
rect 16829 9726 16897 9760
rect 16987 9726 17055 9760
rect 17145 9726 17213 9760
rect 17303 9726 17371 9760
rect 17461 9726 17529 9760
rect 17619 9726 17687 9760
rect 17777 9726 17845 9760
rect 17935 9726 18003 9760
rect 18093 9726 18161 9760
rect 18251 9726 18319 9760
rect 18409 9726 18477 9760
rect 18567 9726 18635 9760
rect 18725 9726 18793 9760
rect 18883 9726 18951 9760
rect 19041 9726 19109 9760
rect 19199 9726 19267 9760
rect 19357 9726 19425 9760
rect 19515 9726 19583 9760
rect 19673 9726 19741 9760
rect 19831 9726 19899 9760
rect 19989 9726 20057 9760
rect 16609 7700 16643 9676
rect 16767 7700 16801 9676
rect 16925 7700 16959 9676
rect 17083 7700 17117 9676
rect 17241 7700 17275 9676
rect 17399 7700 17433 9676
rect 17557 7700 17591 9676
rect 17715 7700 17749 9676
rect 17873 7700 17907 9676
rect 18031 7700 18065 9676
rect 18189 7700 18223 9676
rect 18347 7700 18381 9676
rect 18505 7700 18539 9676
rect 18663 7700 18697 9676
rect 18821 7700 18855 9676
rect 18979 7700 19013 9676
rect 19137 7700 19171 9676
rect 19295 7700 19329 9676
rect 19453 7700 19487 9676
rect 19611 7700 19645 9676
rect 19769 7700 19803 9676
rect 19927 7700 19961 9676
rect 20085 7700 20119 9676
rect 16671 7616 16739 7650
rect 16829 7616 16897 7650
rect 16987 7616 17055 7650
rect 17145 7616 17213 7650
rect 17303 7616 17371 7650
rect 17461 7616 17529 7650
rect 17619 7616 17687 7650
rect 17777 7616 17845 7650
rect 17935 7616 18003 7650
rect 18093 7616 18161 7650
rect 18251 7616 18319 7650
rect 18409 7616 18477 7650
rect 18567 7616 18635 7650
rect 18725 7616 18793 7650
rect 18883 7616 18951 7650
rect 19041 7616 19109 7650
rect 19199 7616 19267 7650
rect 19357 7616 19425 7650
rect 19515 7616 19583 7650
rect 19673 7616 19741 7650
rect 19831 7616 19899 7650
rect 19989 7616 20057 7650
rect 20274 7473 20400 10100
rect 16471 7311 20400 7473
rect 16471 7290 16567 7311
rect 16567 7290 16995 7311
rect 16995 7290 17153 7311
rect 17153 7290 17581 7311
rect 17581 7290 17739 7311
rect 17739 7290 18167 7311
rect 18167 7290 20400 7311
rect 14113 6124 14151 6521
rect 14113 2625 14151 3022
rect 14409 6124 14447 6521
rect 14409 2625 14447 3022
rect 14705 6124 14743 6521
rect 14705 2625 14743 3022
rect 15001 6124 15039 6521
rect 15001 2625 15039 3022
rect 15297 6124 15335 6521
rect 15297 2625 15335 3022
rect 15593 6124 15631 6521
rect 15593 2625 15631 3022
rect 15889 6124 15927 6521
rect 15889 2625 15927 3022
rect 16185 6124 16223 6521
rect 16185 2625 16223 3022
rect 16693 7143 16869 7177
rect 16609 5147 16643 7115
rect 16919 5147 16953 7115
rect 16693 5085 16869 5119
rect 17279 7143 17455 7177
rect 17195 5147 17229 7115
rect 17505 5147 17539 7115
rect 17279 5085 17455 5119
rect 17865 7143 18041 7177
rect 17781 5147 17815 7115
rect 18091 5147 18125 7115
rect 17865 5085 18041 5119
rect 18519 6378 19526 6561
rect 16693 4681 16869 4715
rect 16609 2685 16643 4653
rect 16919 2685 16953 4653
rect 16693 2623 16869 2657
rect 17279 4681 17455 4715
rect 17195 2685 17229 4653
rect 17505 2685 17539 4653
rect 17279 2623 17455 2657
rect 17865 4681 18041 4715
rect 17781 2685 17815 4653
rect 18091 2685 18125 4653
rect 17865 2623 18041 2657
rect 18730 5824 18768 6221
rect 18730 2625 18768 3022
rect 19026 5824 19064 6221
rect 19026 2625 19064 3022
rect 19322 5824 19360 6221
rect 19322 2625 19360 3022
rect 19618 5824 19656 6221
rect 19618 2625 19656 3022
rect 20160 2391 20400 7290
rect 13753 2259 20400 2391
rect 20160 2254 20400 2259
rect 21325 8145 24025 8161
rect 21195 8129 24025 8145
rect 21195 8079 24090 8129
rect 21195 8045 21623 8079
rect 21623 8045 23851 8079
rect 23851 8045 24090 8079
rect 21195 8031 24090 8045
rect 21195 5964 21504 8031
rect 21749 7911 23725 7945
rect 21665 6115 21699 7883
rect 23775 6115 23809 7883
rect 21749 6053 23725 6087
rect 23911 7983 24090 8031
rect 23911 6015 23913 7983
rect 23913 6015 23947 7983
rect 23947 6015 24090 7983
rect 21195 5953 23723 5964
rect 21195 5919 21623 5953
rect 21623 5919 23723 5953
rect 21195 5829 23723 5919
rect 21195 5795 21623 5829
rect 21623 5795 23723 5829
rect 21195 3591 21504 5795
rect 21749 5661 23725 5695
rect 21665 3865 21699 5633
rect 23775 3865 23809 5633
rect 23911 5733 24090 6015
rect 23911 4060 23913 5733
rect 23913 4060 23947 5733
rect 23947 4311 24090 5733
rect 24363 8159 25879 8168
rect 24363 8149 26789 8159
rect 24363 8079 26835 8149
rect 24363 8045 24708 8079
rect 24708 8045 25754 8079
rect 25754 8045 26835 8079
rect 24363 8040 26835 8045
rect 24363 7983 24619 8040
rect 24363 7835 24612 7983
rect 24612 7835 24619 7983
rect 24364 7615 24612 7835
rect 24612 7615 24618 7835
rect 25836 7983 26835 8040
rect 24843 7911 25619 7945
rect 24750 7715 24784 7883
rect 25678 7715 25712 7883
rect 24843 7653 25619 7687
rect 24364 7277 24618 7615
rect 25836 7615 25850 7983
rect 25850 7615 26835 7983
rect 25836 7537 26835 7615
rect 24883 7519 25754 7537
rect 25754 7519 26835 7537
rect 24883 7373 26835 7519
rect 24883 7369 26654 7373
rect 26654 7369 26835 7373
rect 24883 7354 25918 7369
rect 24364 5103 24612 7277
rect 24612 5103 24618 7277
rect 24843 7205 26519 7239
rect 24750 7009 24784 7177
rect 26578 7009 26612 7177
rect 24843 6947 26519 6981
rect 24750 6751 24784 6919
rect 26578 6751 26612 6919
rect 24843 6689 26519 6723
rect 24750 6493 24784 6661
rect 26578 6493 26612 6661
rect 24843 6431 26519 6465
rect 24750 6235 24784 6403
rect 26578 6235 26612 6403
rect 24843 6173 26519 6207
rect 24750 5977 24784 6145
rect 26578 5977 26612 6145
rect 24843 5915 26519 5949
rect 24750 5719 24784 5887
rect 26578 5719 26612 5887
rect 24843 5657 26519 5691
rect 24750 5461 24784 5629
rect 26578 5461 26612 5629
rect 24843 5399 26519 5433
rect 24750 5203 24784 5371
rect 26578 5203 26612 5371
rect 24843 5141 26519 5175
rect 24364 5025 24618 5103
rect 26708 7277 26835 7369
rect 26708 5103 26716 7277
rect 26716 5103 26750 7277
rect 26750 5103 26835 7277
rect 26708 5025 26835 5103
rect 24358 5007 24708 5025
rect 24708 5007 26654 5025
rect 26654 5007 26835 5025
rect 24358 4469 26835 5007
rect 23947 4060 26905 4311
rect 21749 3803 23725 3837
rect 24020 4050 26905 4060
rect 23911 3591 24090 3744
rect 21195 3233 24301 3591
rect 21199 3201 24301 3233
rect 21199 3147 24290 3201
rect 21199 3137 24295 3147
rect 21199 3106 21408 3137
rect 21408 3106 24098 3137
rect 24098 3106 24295 3137
rect 21199 3041 21328 3106
rect 21199 1813 21312 3041
rect 21312 1813 21328 3041
rect 24187 3041 24295 3106
rect 21508 2965 21676 2999
rect 21766 2965 21934 2999
rect 22024 2965 22192 2999
rect 22282 2965 22450 2999
rect 22540 2965 22708 2999
rect 22798 2965 22966 2999
rect 23056 2965 23224 2999
rect 23314 2965 23482 2999
rect 23572 2965 23740 2999
rect 23830 2965 23998 2999
rect 21446 1939 21480 2915
rect 21704 1939 21738 2915
rect 21962 1939 21996 2915
rect 22220 1939 22254 2915
rect 22478 1939 22512 2915
rect 22736 1939 22770 2915
rect 22994 1939 23028 2915
rect 23252 1939 23286 2915
rect 23510 1939 23544 2915
rect 23768 1939 23802 2915
rect 24026 1939 24060 2915
rect 21508 1855 21676 1889
rect 21766 1855 21934 1889
rect 22024 1855 22192 1889
rect 22282 1855 22450 1889
rect 22540 1855 22708 1889
rect 22798 1855 22966 1889
rect 23056 1855 23224 1889
rect 23314 1855 23482 1889
rect 23572 1855 23740 1889
rect 23830 1855 23998 1889
rect 21199 1784 21328 1813
rect 24187 1813 24194 3041
rect 24194 1854 24295 3041
rect 24678 3803 26654 3837
rect 24594 2007 24628 3775
rect 26704 2007 26738 3775
rect 24678 1945 26654 1979
rect 26830 3875 26905 4050
rect 26830 1907 26842 3875
rect 26842 1907 26876 3875
rect 26876 1907 26905 3875
rect 26830 1854 26905 1907
rect 24194 1845 26899 1854
rect 24194 1813 24552 1845
rect 24187 1811 24552 1813
rect 24552 1811 26780 1845
rect 26780 1811 26899 1845
rect 24187 1784 26899 1811
rect 21199 1751 26899 1784
rect 21199 1717 21408 1751
rect 21408 1717 24098 1751
rect 24098 1717 26899 1751
rect 21199 1663 26899 1717
rect 21199 1656 24295 1663
<< metal1 >>
rect 2425 42584 2687 42589
rect 2425 42578 5841 42584
rect 2423 42577 2433 42578
rect 2423 30250 2431 42577
rect 5829 42347 5841 42578
rect 2688 42341 5603 42347
rect 2688 30251 2698 42341
rect 2796 42220 3142 42232
rect 2796 41823 2802 42220
rect 2840 42167 3098 42220
rect 2840 41823 2846 42167
rect 2796 41811 2846 41823
rect 3092 41823 3098 42167
rect 3136 41823 3142 42220
rect 3092 41811 3142 41823
rect 3388 42220 3734 42232
rect 3388 41823 3394 42220
rect 3432 42167 3690 42220
rect 3432 41823 3438 42167
rect 3388 41811 3438 41823
rect 3684 41823 3690 42167
rect 3728 41823 3734 42220
rect 3684 41811 3734 41823
rect 3980 42220 4326 42232
rect 3980 41823 3986 42220
rect 4024 42167 4282 42220
rect 4024 41823 4030 42167
rect 3980 41811 4030 41823
rect 4276 41823 4282 42167
rect 4320 41823 4326 42220
rect 4276 41811 4326 41823
rect 4572 42220 4918 42232
rect 4572 41823 4578 42220
rect 4616 42167 4874 42220
rect 4616 41823 4622 42167
rect 4572 41811 4622 41823
rect 4868 41823 4874 42167
rect 4912 41823 4918 42220
rect 4868 41811 4918 41823
rect 5164 42220 5510 42232
rect 5164 41823 5170 42220
rect 5208 42167 5466 42220
rect 5208 41823 5214 42167
rect 5164 41811 5214 41823
rect 5460 41823 5466 42167
rect 5504 41823 5510 42220
rect 5460 41811 5510 41823
rect 2796 36821 2846 36833
rect 2796 36424 2802 36821
rect 2840 36424 2846 36821
rect 2796 36162 2846 36424
rect 2796 35765 2802 36162
rect 2840 35765 2846 36162
rect 2796 35753 2846 35765
rect 3092 36821 3142 36833
rect 3092 36424 3098 36821
rect 3136 36424 3142 36821
rect 3092 36162 3142 36424
rect 3092 35765 3098 36162
rect 3136 35765 3142 36162
rect 3092 35753 3142 35765
rect 3388 36821 3438 36833
rect 3388 36424 3394 36821
rect 3432 36424 3438 36821
rect 3388 36162 3438 36424
rect 3388 35765 3394 36162
rect 3432 35765 3438 36162
rect 3388 35753 3438 35765
rect 3684 36821 3734 36833
rect 3684 36424 3690 36821
rect 3728 36424 3734 36821
rect 3684 36162 3734 36424
rect 3684 35765 3690 36162
rect 3728 35765 3734 36162
rect 3684 35753 3734 35765
rect 3980 36821 4030 36833
rect 3980 36424 3986 36821
rect 4024 36424 4030 36821
rect 3980 36162 4030 36424
rect 3980 35765 3986 36162
rect 4024 35765 4030 36162
rect 3980 35753 4030 35765
rect 4276 36821 4326 36833
rect 4276 36424 4282 36821
rect 4320 36424 4326 36821
rect 4276 36162 4326 36424
rect 4276 35765 4282 36162
rect 4320 35765 4326 36162
rect 4276 35753 4326 35765
rect 4572 36821 4622 36833
rect 4572 36424 4578 36821
rect 4616 36424 4622 36821
rect 4572 36162 4622 36424
rect 4572 35765 4578 36162
rect 4616 35765 4622 36162
rect 4572 35753 4622 35765
rect 4868 36821 4918 36833
rect 4868 36424 4874 36821
rect 4912 36424 4918 36821
rect 4868 36162 4918 36424
rect 4868 35765 4874 36162
rect 4912 35765 4918 36162
rect 4868 35753 4918 35765
rect 5164 36821 5214 36833
rect 5164 36424 5170 36821
rect 5208 36424 5214 36821
rect 5164 36162 5214 36424
rect 5164 35765 5170 36162
rect 5208 35765 5214 36162
rect 5164 35753 5214 35765
rect 5460 36821 5510 36833
rect 5460 36424 5466 36821
rect 5504 36424 5510 36821
rect 5460 36162 5510 36424
rect 5460 35765 5466 36162
rect 5504 35765 5510 36162
rect 5460 35753 5510 35765
rect 5593 31000 5603 42341
rect 5815 42341 5841 42347
rect 5815 31000 5825 42341
rect 6020 31303 10895 31309
rect 6020 31147 6032 31303
rect 6020 31112 6028 31147
rect 10883 31118 10895 31303
rect 2796 30766 2846 30775
rect 2774 30366 2784 30766
rect 2856 30366 2866 30766
rect 3092 30763 3142 30775
rect 3092 30366 3098 30763
rect 3136 30419 3142 30763
rect 3388 30763 3438 30775
rect 3388 30419 3394 30763
rect 3136 30366 3394 30419
rect 3432 30366 3438 30763
rect 2796 30354 2846 30366
rect 3092 30354 3438 30366
rect 3684 30763 3734 30775
rect 3684 30366 3690 30763
rect 3728 30419 3734 30763
rect 3980 30763 4030 30775
rect 3980 30419 3986 30763
rect 3728 30366 3986 30419
rect 4024 30366 4030 30763
rect 3684 30354 4030 30366
rect 4276 30763 4326 30775
rect 4276 30366 4282 30763
rect 4320 30419 4326 30763
rect 4572 30763 4622 30775
rect 4572 30419 4578 30763
rect 4320 30366 4578 30419
rect 4616 30366 4622 30763
rect 4276 30354 4622 30366
rect 4868 30763 4918 30775
rect 4868 30366 4874 30763
rect 4912 30419 4918 30763
rect 5164 30763 5214 30775
rect 5460 30763 5510 30775
rect 5164 30419 5170 30763
rect 4912 30366 5170 30419
rect 5208 30366 5214 30763
rect 5449 30366 5459 30763
rect 5511 30366 5521 30763
rect 4868 30354 5214 30366
rect 5460 30354 5510 30366
rect 5607 30251 5613 31000
rect 2688 30250 5613 30251
rect 5815 30251 5821 31000
rect 6022 30542 6028 31112
rect 6019 30450 6028 30542
rect 6143 31112 10759 31118
rect 6143 30542 6149 31112
rect 6283 30999 8275 31005
rect 6283 30965 6295 30999
rect 8263 30965 8275 30999
rect 6283 30959 8275 30965
rect 8609 30999 10601 31005
rect 8609 30965 8621 30999
rect 10589 30965 10601 30999
rect 8609 30959 10601 30965
rect 6227 30906 6273 30918
rect 6227 30830 6233 30906
rect 6267 30830 6273 30906
rect 8285 30906 8331 30918
rect 6214 30730 6224 30830
rect 6276 30730 6286 30830
rect 8285 30730 8291 30906
rect 8325 30784 8331 30906
rect 8553 30906 8599 30918
rect 10611 30906 10657 30918
rect 8553 30784 8559 30906
rect 8325 30730 8559 30784
rect 8593 30730 8599 30906
rect 10592 30806 10602 30906
rect 10666 30806 10676 30906
rect 6227 30718 6273 30730
rect 8285 30718 8599 30730
rect 10611 30730 10617 30806
rect 10651 30730 10657 30806
rect 10611 30718 10657 30730
rect 6285 30677 6295 30679
rect 6283 30631 6295 30677
rect 6548 30677 6558 30679
rect 10219 30677 10229 30686
rect 6548 30671 10229 30677
rect 10589 30677 10599 30686
rect 8263 30637 8621 30671
rect 6285 30622 6295 30631
rect 6548 30631 10229 30637
rect 6548 30622 6558 30631
rect 10219 30613 10229 30631
rect 10589 30631 10601 30677
rect 10589 30613 10599 30631
rect 10749 30542 10759 31112
rect 6143 30536 10759 30542
rect 10874 31112 10895 31118
rect 10874 30542 10884 31112
rect 10874 30536 10894 30542
rect 6019 30351 6031 30450
rect 10882 30351 10894 30536
rect 6019 30345 10894 30351
rect 2419 30063 2429 30250
rect 2425 30058 2491 30063
rect 5815 30058 5827 30251
rect 2425 30052 5827 30058
rect 2425 30051 2687 30052
rect 7365 28349 7496 28352
rect 17595 28349 17794 28352
rect 7358 28343 17794 28349
rect 7358 28190 7370 28343
rect 17591 28190 17794 28343
rect 7358 28184 7371 28190
rect 7365 27985 7371 28184
rect 7104 27983 7371 27985
rect 6226 27582 6236 27983
rect 7095 27582 7371 27983
rect 5736 24621 5987 24633
rect 5732 19960 5742 24621
rect 5981 24620 5991 24621
rect 7365 24620 7371 27582
rect 5981 24614 7371 24620
rect 7490 28184 13405 28190
rect 7490 28103 7496 28184
rect 13399 28103 13405 28184
rect 7490 28097 8013 28103
rect 7490 28059 7604 28097
rect 8001 28059 8013 28097
rect 7490 28053 8013 28059
rect 9891 28097 13405 28103
rect 9891 28059 9903 28097
rect 10300 28059 10562 28097
rect 10959 28059 12861 28097
rect 13258 28059 13405 28097
rect 9891 28053 13405 28059
rect 7490 24857 7496 28053
rect 12851 27807 12861 27808
rect 7592 27801 8013 27807
rect 7592 27763 7604 27801
rect 8001 27763 8013 27801
rect 7592 27757 8013 27763
rect 9891 27801 10971 27807
rect 9891 27763 9903 27801
rect 10300 27763 10562 27801
rect 10959 27763 10971 27801
rect 9891 27757 10971 27763
rect 12849 27757 12861 27807
rect 13258 27807 13268 27808
rect 7592 27511 7674 27757
rect 12851 27756 12861 27757
rect 13258 27757 13270 27807
rect 13258 27756 13268 27757
rect 7592 27505 8013 27511
rect 7592 27467 7604 27505
rect 8001 27467 8013 27505
rect 7592 27461 8013 27467
rect 9891 27505 10971 27511
rect 9891 27467 9903 27505
rect 10300 27467 10562 27505
rect 10959 27467 10971 27505
rect 9891 27461 10971 27467
rect 12849 27505 13270 27511
rect 12849 27467 12861 27505
rect 13258 27467 13270 27505
rect 12849 27461 13270 27467
rect 13188 27215 13270 27461
rect 7592 27209 8013 27215
rect 7592 27171 7604 27209
rect 8001 27171 8013 27209
rect 7592 27165 8013 27171
rect 9891 27209 10971 27215
rect 9891 27171 9903 27209
rect 10300 27171 10562 27209
rect 10959 27171 10971 27209
rect 9891 27165 10971 27171
rect 12849 27209 13270 27215
rect 12849 27171 12861 27209
rect 13258 27171 13270 27209
rect 12849 27165 13270 27171
rect 7592 26919 7674 27165
rect 7592 26913 8013 26919
rect 7592 26875 7604 26913
rect 8001 26875 8013 26913
rect 7592 26869 8013 26875
rect 9891 26913 10971 26919
rect 9891 26875 9903 26913
rect 10300 26875 10562 26913
rect 10959 26875 10971 26913
rect 9891 26869 10971 26875
rect 12849 26913 13270 26919
rect 12849 26875 12861 26913
rect 13258 26875 13270 26913
rect 12849 26869 13270 26875
rect 13188 26623 13270 26869
rect 7592 26617 8013 26623
rect 7592 26579 7604 26617
rect 8001 26579 8013 26617
rect 7592 26573 8013 26579
rect 9891 26617 10971 26623
rect 9891 26579 9903 26617
rect 10300 26579 10562 26617
rect 10959 26579 10971 26617
rect 9891 26573 10971 26579
rect 12849 26617 13270 26623
rect 12849 26579 12861 26617
rect 13258 26579 13270 26617
rect 12849 26573 13270 26579
rect 7592 26327 7674 26573
rect 7592 26321 8013 26327
rect 7592 26283 7604 26321
rect 8001 26283 8013 26321
rect 7592 26277 8013 26283
rect 9891 26321 10971 26327
rect 9891 26283 9903 26321
rect 10300 26283 10562 26321
rect 10959 26283 10971 26321
rect 9891 26277 10971 26283
rect 12849 26321 13270 26327
rect 12849 26283 12861 26321
rect 13258 26283 13270 26321
rect 12849 26277 13270 26283
rect 13188 26031 13270 26277
rect 7592 26025 8013 26031
rect 7592 25987 7604 26025
rect 8001 25987 8013 26025
rect 7592 25981 8013 25987
rect 9891 26025 10971 26031
rect 9891 25987 9903 26025
rect 10300 25987 10562 26025
rect 10959 25987 10971 26025
rect 9891 25981 10971 25987
rect 12849 26025 13270 26031
rect 12849 25987 12861 26025
rect 13258 25987 13270 26025
rect 12849 25981 13270 25987
rect 7592 25735 7674 25981
rect 7592 25729 8013 25735
rect 7592 25691 7604 25729
rect 8001 25691 8013 25729
rect 7592 25685 8013 25691
rect 9891 25729 10971 25735
rect 9891 25691 9903 25729
rect 10300 25691 10562 25729
rect 10959 25691 10971 25729
rect 9891 25685 10971 25691
rect 12849 25729 13270 25735
rect 12849 25691 12861 25729
rect 13258 25691 13270 25729
rect 12849 25685 13270 25691
rect 13188 25439 13270 25685
rect 7592 25433 8013 25439
rect 7592 25395 7604 25433
rect 8001 25395 8013 25433
rect 7592 25389 8013 25395
rect 9891 25433 10971 25439
rect 9891 25395 9903 25433
rect 10300 25395 10562 25433
rect 10959 25395 10971 25433
rect 9891 25389 10971 25395
rect 12849 25433 13270 25439
rect 12849 25395 12861 25433
rect 13258 25395 13270 25433
rect 12849 25389 13270 25395
rect 7592 25143 7674 25389
rect 12948 25143 12958 25144
rect 7592 25137 8013 25143
rect 7592 25099 7604 25137
rect 8001 25099 8013 25137
rect 7592 25093 8013 25099
rect 9891 25137 10971 25143
rect 9891 25099 9903 25137
rect 10300 25099 10562 25137
rect 10959 25099 10971 25137
rect 9891 25093 10971 25099
rect 12849 25137 12958 25143
rect 13258 25143 13268 25144
rect 12849 25099 12861 25137
rect 12849 25093 12958 25099
rect 12948 25092 12958 25093
rect 13258 25093 13270 25143
rect 13258 25092 13268 25093
rect 7490 24847 7612 24857
rect 13399 24848 13405 28053
rect 17590 28168 17794 28190
rect 13844 28044 14739 28050
rect 13844 27184 13850 28044
rect 13986 27892 14596 27923
rect 13986 27858 14031 27892
rect 14065 27858 14131 27892
rect 14165 27858 14231 27892
rect 14265 27858 14331 27892
rect 14365 27858 14431 27892
rect 14465 27858 14531 27892
rect 14565 27858 14596 27892
rect 13986 27818 14596 27858
rect 14727 27825 14739 28044
rect 15181 28044 16084 28050
rect 15181 27825 15193 28044
rect 14727 27819 15193 27825
rect 15330 27892 15940 27923
rect 15330 27858 15375 27892
rect 15409 27858 15475 27892
rect 15509 27858 15575 27892
rect 15609 27858 15675 27892
rect 15709 27858 15775 27892
rect 15809 27858 15875 27892
rect 15909 27858 15940 27892
rect 13976 27344 13986 27818
rect 14066 27792 14596 27818
rect 14066 27758 14131 27792
rect 14165 27758 14231 27792
rect 14265 27758 14331 27792
rect 14365 27758 14431 27792
rect 14465 27758 14531 27792
rect 14565 27758 14596 27792
rect 14066 27750 14596 27758
rect 15330 27792 15940 27858
rect 16072 27814 16084 28044
rect 16526 28044 17424 28050
rect 16526 27814 16538 28044
rect 16072 27808 16538 27814
rect 16674 27892 17284 27923
rect 16674 27858 16719 27892
rect 16753 27858 16819 27892
rect 16853 27858 16919 27892
rect 16953 27858 17019 27892
rect 17053 27858 17119 27892
rect 17153 27858 17219 27892
rect 17253 27858 17284 27892
rect 15330 27758 15375 27792
rect 15409 27758 15475 27792
rect 15509 27758 15575 27792
rect 15609 27758 15675 27792
rect 15709 27758 15775 27792
rect 15809 27758 15875 27792
rect 15909 27758 15940 27792
rect 15330 27750 15940 27758
rect 14066 27744 15940 27750
rect 16674 27792 17284 27858
rect 16674 27758 16719 27792
rect 16753 27758 16819 27792
rect 16853 27758 16919 27792
rect 16953 27758 17019 27792
rect 17053 27758 17119 27792
rect 17153 27758 17219 27792
rect 17253 27758 17284 27792
rect 16674 27744 17284 27758
rect 14066 27692 17284 27744
rect 14066 27658 14131 27692
rect 14165 27658 14231 27692
rect 14265 27658 14331 27692
rect 14365 27658 14431 27692
rect 14465 27658 14531 27692
rect 14565 27658 15375 27692
rect 15409 27658 15475 27692
rect 15509 27658 15575 27692
rect 15609 27658 15675 27692
rect 15709 27658 15775 27692
rect 15809 27658 15875 27692
rect 15909 27658 16719 27692
rect 16753 27658 16819 27692
rect 16853 27658 16919 27692
rect 16953 27658 17019 27692
rect 17053 27658 17119 27692
rect 17153 27658 17219 27692
rect 17253 27658 17284 27692
rect 14066 27592 17284 27658
rect 14066 27558 14131 27592
rect 14165 27558 14231 27592
rect 14265 27558 14331 27592
rect 14365 27558 14431 27592
rect 14465 27558 14531 27592
rect 14565 27558 15375 27592
rect 15409 27558 15475 27592
rect 15509 27558 15575 27592
rect 15609 27558 15675 27592
rect 15709 27558 15775 27592
rect 15809 27558 15875 27592
rect 15909 27558 16719 27592
rect 16753 27558 16819 27592
rect 16853 27558 16919 27592
rect 16953 27558 17019 27592
rect 17053 27558 17119 27592
rect 17153 27558 17219 27592
rect 17253 27558 17284 27592
rect 14066 27492 17284 27558
rect 14066 27458 14131 27492
rect 14165 27458 14231 27492
rect 14265 27458 14331 27492
rect 14365 27458 14431 27492
rect 14465 27458 14531 27492
rect 14565 27470 15375 27492
rect 14565 27458 14596 27470
rect 14066 27392 14596 27458
rect 14066 27358 14131 27392
rect 14165 27358 14231 27392
rect 14265 27358 14331 27392
rect 14365 27358 14431 27392
rect 14465 27358 14531 27392
rect 14565 27358 14596 27392
rect 15330 27458 15375 27470
rect 15409 27458 15475 27492
rect 15509 27458 15575 27492
rect 15609 27458 15675 27492
rect 15709 27458 15775 27492
rect 15809 27458 15875 27492
rect 15909 27464 16719 27492
rect 15909 27458 15940 27464
rect 15330 27392 15940 27458
rect 14066 27344 14596 27358
rect 13986 27313 14596 27344
rect 14756 27372 15184 27384
rect 13844 27172 14088 27184
rect 14082 26863 14088 27172
rect 13844 26851 14088 26863
rect 13844 25838 13850 26851
rect 14143 26579 14452 27313
rect 14756 27181 14762 27372
rect 14538 27175 14762 27181
rect 15178 27181 15184 27372
rect 15330 27358 15375 27392
rect 15409 27358 15475 27392
rect 15509 27358 15575 27392
rect 15609 27358 15675 27392
rect 15709 27358 15775 27392
rect 15809 27358 15875 27392
rect 15909 27358 15940 27392
rect 16674 27458 16719 27464
rect 16753 27458 16819 27492
rect 16853 27458 16919 27492
rect 16953 27458 17019 27492
rect 17053 27458 17119 27492
rect 17153 27458 17219 27492
rect 17253 27458 17284 27492
rect 16674 27392 17284 27458
rect 15330 27313 15940 27358
rect 16086 27372 16514 27384
rect 16086 27181 16092 27372
rect 15178 27175 16092 27181
rect 16508 27181 16514 27372
rect 16674 27358 16719 27392
rect 16753 27358 16819 27392
rect 16853 27358 16919 27392
rect 16953 27358 17019 27392
rect 17053 27358 17119 27392
rect 17153 27358 17219 27392
rect 17253 27358 17284 27392
rect 16674 27313 17284 27358
rect 16508 27175 16776 27181
rect 14538 26877 14550 27175
rect 16764 26877 16776 27175
rect 14538 26871 14762 26877
rect 13986 26548 14596 26579
rect 13986 26514 14031 26548
rect 14065 26514 14131 26548
rect 14165 26514 14231 26548
rect 14265 26514 14331 26548
rect 14365 26514 14431 26548
rect 14465 26514 14531 26548
rect 14565 26514 14596 26548
rect 13986 26448 14596 26514
rect 13986 26414 14031 26448
rect 14065 26414 14131 26448
rect 14165 26414 14231 26448
rect 14265 26414 14331 26448
rect 14365 26414 14431 26448
rect 14465 26414 14531 26448
rect 14565 26414 14596 26448
rect 13986 26348 14596 26414
rect 13986 26314 14031 26348
rect 14065 26314 14131 26348
rect 14165 26314 14231 26348
rect 14265 26314 14331 26348
rect 14365 26314 14431 26348
rect 14465 26314 14531 26348
rect 14565 26314 14596 26348
rect 13986 26248 14596 26314
rect 13986 26214 14031 26248
rect 14065 26214 14131 26248
rect 14165 26214 14231 26248
rect 14265 26214 14331 26248
rect 14365 26214 14431 26248
rect 14465 26214 14531 26248
rect 14565 26214 14596 26248
rect 13986 26148 14596 26214
rect 13986 26114 14031 26148
rect 14065 26114 14131 26148
rect 14165 26114 14231 26148
rect 14265 26114 14331 26148
rect 14365 26114 14431 26148
rect 14465 26114 14531 26148
rect 14565 26114 14596 26148
rect 13986 26048 14596 26114
rect 13986 26014 14031 26048
rect 14065 26014 14131 26048
rect 14165 26014 14231 26048
rect 14265 26014 14331 26048
rect 14365 26014 14431 26048
rect 14465 26014 14531 26048
rect 14565 26014 14596 26048
rect 13986 25969 14596 26014
rect 13844 25826 14088 25838
rect 14082 25517 14088 25826
rect 13256 24847 13405 24848
rect 7490 24841 13405 24847
rect 7490 24803 7604 24841
rect 8001 24803 9903 24841
rect 10300 24803 10562 24841
rect 10959 24803 12861 24841
rect 13258 24803 13405 24841
rect 7490 24797 13405 24803
rect 7490 24787 7612 24797
rect 7490 24620 7496 24787
rect 7490 24614 11244 24620
rect 11232 24608 11244 24614
rect 13399 24608 13405 24797
rect 11232 24602 13405 24608
rect 13844 25505 14088 25517
rect 13844 24502 13850 25505
rect 14140 25235 14449 25969
rect 14756 25832 14762 26871
rect 14569 25826 14762 25832
rect 15178 26871 16092 26877
rect 15178 25832 15184 26871
rect 15330 26548 15940 26579
rect 15330 26514 15375 26548
rect 15409 26514 15475 26548
rect 15509 26514 15575 26548
rect 15609 26514 15675 26548
rect 15709 26514 15775 26548
rect 15809 26514 15875 26548
rect 15909 26514 15940 26548
rect 15330 26448 15940 26514
rect 15330 26414 15375 26448
rect 15409 26414 15475 26448
rect 15509 26414 15575 26448
rect 15609 26414 15675 26448
rect 15709 26414 15775 26448
rect 15809 26414 15875 26448
rect 15909 26414 15940 26448
rect 15330 26348 15940 26414
rect 15330 26314 15375 26348
rect 15409 26314 15475 26348
rect 15509 26314 15575 26348
rect 15609 26314 15675 26348
rect 15709 26314 15775 26348
rect 15809 26314 15875 26348
rect 15909 26314 15940 26348
rect 15330 26248 15940 26314
rect 15330 26214 15375 26248
rect 15409 26214 15475 26248
rect 15509 26214 15575 26248
rect 15609 26214 15675 26248
rect 15709 26214 15775 26248
rect 15809 26214 15875 26248
rect 15909 26214 15940 26248
rect 15330 26148 15940 26214
rect 15330 26114 15375 26148
rect 15409 26114 15475 26148
rect 15509 26114 15575 26148
rect 15609 26114 15675 26148
rect 15709 26114 15775 26148
rect 15809 26114 15875 26148
rect 15909 26114 15940 26148
rect 15330 26070 15940 26114
rect 15330 26048 15378 26070
rect 15907 26048 15940 26070
rect 15330 26014 15375 26048
rect 15909 26014 15940 26048
rect 15330 25984 15378 26014
rect 15907 25984 15940 26014
rect 15330 25969 15940 25984
rect 16086 25832 16092 26871
rect 15178 25826 16092 25832
rect 16508 26871 16776 26877
rect 16508 25832 16514 26871
rect 16839 26579 17148 27313
rect 17418 27191 17424 28044
rect 17189 27179 17424 27191
rect 17590 28044 17602 28168
rect 17189 26870 17195 27179
rect 17189 26858 17424 26870
rect 16674 26548 17284 26579
rect 16674 26514 16719 26548
rect 16753 26514 16819 26548
rect 16853 26514 16919 26548
rect 16953 26514 17019 26548
rect 17053 26514 17119 26548
rect 17153 26514 17219 26548
rect 17253 26514 17284 26548
rect 16674 26448 17284 26514
rect 16674 26414 16719 26448
rect 16753 26414 16819 26448
rect 16853 26414 16919 26448
rect 16953 26414 17019 26448
rect 17053 26414 17119 26448
rect 17153 26414 17219 26448
rect 17253 26414 17284 26448
rect 16674 26348 17284 26414
rect 16674 26314 16719 26348
rect 16753 26314 16819 26348
rect 16853 26314 16919 26348
rect 16953 26314 17019 26348
rect 17053 26314 17119 26348
rect 17153 26314 17219 26348
rect 17253 26314 17284 26348
rect 16674 26248 17284 26314
rect 16674 26214 16719 26248
rect 16753 26214 16819 26248
rect 16853 26214 16919 26248
rect 16953 26214 17019 26248
rect 17053 26214 17119 26248
rect 17153 26214 17219 26248
rect 17253 26214 17284 26248
rect 16674 26148 17284 26214
rect 16674 26114 16719 26148
rect 16753 26114 16819 26148
rect 16853 26114 16919 26148
rect 16953 26114 17019 26148
rect 17053 26114 17119 26148
rect 17153 26114 17219 26148
rect 17253 26114 17284 26148
rect 16674 26048 17284 26114
rect 16674 26014 16719 26048
rect 16753 26014 16819 26048
rect 16853 26014 16919 26048
rect 16953 26014 17019 26048
rect 17053 26014 17119 26048
rect 17153 26014 17219 26048
rect 17253 26014 17284 26048
rect 16674 25969 17284 26014
rect 16508 25826 16765 25832
rect 14569 25520 14581 25826
rect 16753 25520 16765 25826
rect 14569 25514 14762 25520
rect 13986 25204 14596 25235
rect 13986 25170 14031 25204
rect 14065 25170 14131 25204
rect 14165 25170 14231 25204
rect 14265 25170 14331 25204
rect 14365 25170 14431 25204
rect 14465 25170 14531 25204
rect 14565 25170 14596 25204
rect 13986 25104 14596 25170
rect 13986 25070 14031 25104
rect 14065 25070 14131 25104
rect 14165 25070 14231 25104
rect 14265 25070 14331 25104
rect 14365 25070 14431 25104
rect 14465 25070 14531 25104
rect 14565 25070 14596 25104
rect 14756 25105 14762 25514
rect 15178 25514 16092 25520
rect 15178 25105 15184 25514
rect 14756 25093 15184 25105
rect 15330 25204 15940 25235
rect 15330 25170 15375 25204
rect 15409 25170 15475 25204
rect 15509 25170 15575 25204
rect 15609 25170 15675 25204
rect 15709 25170 15775 25204
rect 15809 25170 15875 25204
rect 15909 25170 15940 25204
rect 15330 25104 15940 25170
rect 13986 25050 14596 25070
rect 15330 25070 15375 25104
rect 15409 25070 15475 25104
rect 15509 25070 15575 25104
rect 15609 25070 15675 25104
rect 15709 25070 15775 25104
rect 15809 25070 15875 25104
rect 15909 25070 15940 25104
rect 16086 25105 16092 25514
rect 16508 25514 16765 25520
rect 16508 25105 16514 25514
rect 16844 25235 17153 25969
rect 17418 25857 17424 26858
rect 17204 25845 17424 25857
rect 17204 25501 17210 25845
rect 17204 25489 17424 25501
rect 16086 25093 16514 25105
rect 16674 25204 17284 25235
rect 16674 25170 16719 25204
rect 16753 25170 16819 25204
rect 16853 25170 16919 25204
rect 16953 25170 17019 25204
rect 17053 25170 17119 25204
rect 17153 25170 17219 25204
rect 17253 25170 17284 25204
rect 16674 25104 17284 25170
rect 15330 25050 15940 25070
rect 13986 25047 15940 25050
rect 16674 25070 16719 25104
rect 16753 25070 16819 25104
rect 16853 25070 16919 25104
rect 16953 25070 17019 25104
rect 17053 25070 17119 25104
rect 17153 25070 17219 25104
rect 17253 25070 17284 25104
rect 16674 25047 17284 25070
rect 13986 25004 17284 25047
rect 13986 24970 14031 25004
rect 14065 24970 14131 25004
rect 14165 24970 14231 25004
rect 14265 24970 14331 25004
rect 14365 24970 14431 25004
rect 14465 24970 14531 25004
rect 14565 24970 15375 25004
rect 15409 24970 15475 25004
rect 15509 24970 15575 25004
rect 15609 24970 15675 25004
rect 15709 24970 15775 25004
rect 15809 24970 15875 25004
rect 15909 24970 16719 25004
rect 16753 24970 16819 25004
rect 16853 24970 16919 25004
rect 16953 24970 17019 25004
rect 17053 24970 17119 25004
rect 17153 24970 17219 25004
rect 17253 24970 17284 25004
rect 13986 24904 17284 24970
rect 13986 24870 14031 24904
rect 14065 24870 14131 24904
rect 14165 24870 14231 24904
rect 14265 24870 14331 24904
rect 14365 24870 14431 24904
rect 14465 24870 14531 24904
rect 14565 24870 15375 24904
rect 15409 24870 15475 24904
rect 15509 24870 15575 24904
rect 15609 24870 15675 24904
rect 15709 24870 15775 24904
rect 15809 24870 15875 24904
rect 15909 24870 16719 24904
rect 16753 24870 16819 24904
rect 16853 24870 16919 24904
rect 16953 24870 17019 24904
rect 17053 24870 17119 24904
rect 17153 24870 17219 24904
rect 17253 24870 17284 24904
rect 13986 24804 17284 24870
rect 13986 24770 14031 24804
rect 14065 24770 14131 24804
rect 14165 24770 14231 24804
rect 14265 24770 14331 24804
rect 14365 24770 14431 24804
rect 14465 24770 14531 24804
rect 14565 24770 15375 24804
rect 15409 24770 15475 24804
rect 15509 24770 15575 24804
rect 15609 24770 15675 24804
rect 15709 24770 15775 24804
rect 15809 24770 15875 24804
rect 15909 24770 16719 24804
rect 16753 24770 16819 24804
rect 16853 24770 16919 24804
rect 16953 24770 17019 24804
rect 17053 24770 17119 24804
rect 17153 24770 17219 24804
rect 17253 24770 17284 24804
rect 13986 24704 14596 24770
rect 15330 24767 17284 24770
rect 13986 24670 14031 24704
rect 14065 24670 14131 24704
rect 14165 24670 14231 24704
rect 14265 24670 14331 24704
rect 14365 24670 14431 24704
rect 14465 24670 14531 24704
rect 14565 24670 14596 24704
rect 13986 24625 14596 24670
rect 14731 24716 15197 24722
rect 14731 24502 14743 24716
rect 13844 24496 14743 24502
rect 15185 24502 15197 24716
rect 15330 24704 15940 24767
rect 15330 24670 15375 24704
rect 15409 24670 15475 24704
rect 15509 24670 15575 24704
rect 15609 24670 15675 24704
rect 15709 24670 15775 24704
rect 15809 24670 15875 24704
rect 15909 24670 15940 24704
rect 15330 24625 15940 24670
rect 16076 24712 16542 24718
rect 16076 24502 16088 24712
rect 15185 24496 16088 24502
rect 16530 24502 16542 24712
rect 16674 24704 17284 24767
rect 16674 24670 16719 24704
rect 16753 24670 16819 24704
rect 16853 24670 16919 24704
rect 16953 24670 17019 24704
rect 17053 24670 17119 24704
rect 17153 24670 17219 24704
rect 17253 24670 17284 24704
rect 16674 24625 17284 24670
rect 17418 24502 17424 25489
rect 16530 24496 17424 24502
rect 17590 24502 17596 28044
rect 17590 24496 17604 24502
rect 17592 24393 17604 24496
rect 17592 24387 17610 24393
rect 12844 24205 13517 24211
rect 12844 24204 12854 24205
rect 13505 24204 13517 24205
rect 11232 24198 11244 24204
rect 13505 24198 15561 24204
rect 5730 19731 5742 19960
rect 5981 24192 6428 24198
rect 5981 19960 5991 24192
rect 6152 24102 6252 24108
rect 6148 24068 6164 24102
rect 6240 24068 6256 24102
rect 6152 24062 6180 24068
rect 6074 24040 6120 24057
rect 6170 24050 6180 24062
rect 6240 24062 6252 24068
rect 6240 24050 6250 24062
rect 6074 20072 6080 24040
rect 6114 23774 6120 24040
rect 6284 24040 6330 24056
rect 6284 23961 6290 24040
rect 6324 23961 6330 24040
rect 6270 23774 6280 23961
rect 6114 22961 6280 23774
rect 6332 22961 6342 23961
rect 6114 20332 6290 22961
rect 6114 20072 6120 20332
rect 6074 20044 6120 20072
rect 6284 20072 6290 20332
rect 6324 20072 6330 22961
rect 6152 20044 6180 20050
rect 6240 20044 6252 20050
rect 6284 20044 6330 20072
rect 6074 20010 6164 20044
rect 6240 20010 6330 20044
rect 6152 20004 6180 20010
rect 6170 19998 6180 20004
rect 6240 20004 6252 20010
rect 6240 19998 6250 20004
rect 6422 19960 6428 24192
rect 5981 19954 6428 19960
rect 6462 24192 6914 24198
rect 6462 19960 6468 24192
rect 6638 24102 6738 24108
rect 6638 24062 6650 24102
rect 6726 24068 6738 24102
rect 6560 24040 6606 24052
rect 6640 24050 6650 24062
rect 6710 24062 6738 24068
rect 6710 24050 6720 24062
rect 6560 23961 6566 24040
rect 6600 23961 6606 24040
rect 6770 24040 6816 24052
rect 6770 23961 6776 24040
rect 6810 23961 6816 24040
rect 6548 22961 6558 23961
rect 6610 23774 6620 23961
rect 6758 23774 6768 23961
rect 6610 22961 6768 23774
rect 6820 22961 6830 23961
rect 6560 20072 6566 22961
rect 6600 20332 6776 22961
rect 6600 20072 6606 20332
rect 6560 20060 6606 20072
rect 6770 20072 6776 20332
rect 6810 20072 6816 22961
rect 6770 20060 6816 20072
rect 6638 20044 6738 20050
rect 6638 20010 6650 20044
rect 6638 20004 6666 20010
rect 6656 19992 6666 20004
rect 6726 20004 6738 20044
rect 6726 19992 6736 20004
rect 6908 19960 6914 24192
rect 6462 19954 6914 19960
rect 6948 24192 7400 24198
rect 6948 19960 6954 24192
rect 7142 24108 7152 24120
rect 7124 24102 7152 24108
rect 7212 24108 7222 24120
rect 7124 24068 7136 24102
rect 7212 24068 7224 24108
rect 7124 24062 7224 24068
rect 7046 24040 7092 24052
rect 7046 23963 7052 24040
rect 7086 23963 7092 24040
rect 7256 24040 7302 24052
rect 7036 22963 7046 23963
rect 7098 23774 7108 23963
rect 7256 23774 7262 24040
rect 7098 22963 7262 23774
rect 7046 20072 7052 22963
rect 7086 20332 7262 22963
rect 7086 20072 7092 20332
rect 7046 20060 7092 20072
rect 7256 20072 7262 20332
rect 7296 20072 7302 24040
rect 7256 20060 7302 20072
rect 7124 20044 7224 20050
rect 7124 20004 7136 20044
rect 7212 20010 7224 20044
rect 7126 19992 7136 20004
rect 7196 20004 7224 20010
rect 7196 19992 7206 20004
rect 7394 19960 7400 24192
rect 6948 19954 7400 19960
rect 7434 24192 7886 24198
rect 7434 19960 7440 24192
rect 7628 24108 7638 24120
rect 7610 24102 7638 24108
rect 7698 24108 7708 24120
rect 7698 24102 7710 24108
rect 7610 24068 7622 24102
rect 7698 24068 7714 24102
rect 7610 24062 7710 24068
rect 7532 24040 7578 24056
rect 7532 20072 7538 24040
rect 7572 23783 7578 24040
rect 7742 24040 7788 24058
rect 7742 23966 7748 24040
rect 7782 23966 7788 24040
rect 7727 23783 7737 23966
rect 7572 22966 7737 23783
rect 7789 22966 7799 23966
rect 7572 20337 7748 22966
rect 7572 20072 7578 20337
rect 7532 20044 7578 20072
rect 7742 20072 7748 20337
rect 7782 20072 7788 22966
rect 7610 20044 7710 20050
rect 7742 20044 7788 20072
rect 7532 20010 7622 20044
rect 7698 20010 7788 20044
rect 7610 20004 7622 20010
rect 7612 19992 7622 20004
rect 7682 20009 7788 20010
rect 7682 20004 7710 20009
rect 7682 19992 7692 20004
rect 7880 19960 7886 24192
rect 7434 19954 7886 19960
rect 7920 24192 8372 24198
rect 7920 19960 7926 24192
rect 8098 24108 8108 24120
rect 8096 24068 8108 24108
rect 8168 24108 8178 24120
rect 8168 24102 8196 24108
rect 8184 24068 8196 24102
rect 8096 24062 8196 24068
rect 8018 24040 8064 24052
rect 8018 23966 8024 24040
rect 8058 23966 8064 24040
rect 8228 24040 8274 24052
rect 8006 22966 8016 23966
rect 8068 23783 8078 23966
rect 8228 23964 8234 24040
rect 8268 23964 8274 24040
rect 8215 23783 8225 23964
rect 8068 22966 8225 23783
rect 8018 20072 8024 22966
rect 8058 22964 8225 22966
rect 8277 22964 8287 23964
rect 8058 20337 8234 22964
rect 8058 20072 8064 20337
rect 8018 20060 8064 20072
rect 8228 20072 8234 20337
rect 8268 20072 8274 22964
rect 8228 20060 8274 20072
rect 8096 20044 8196 20050
rect 8096 20010 8108 20044
rect 8096 20004 8124 20010
rect 8114 19992 8124 20004
rect 8184 20004 8196 20044
rect 8184 19992 8194 20004
rect 8366 19960 8372 24192
rect 7920 19954 8372 19960
rect 8406 24192 8858 24198
rect 8406 19960 8412 24192
rect 8600 24108 8610 24120
rect 8582 24102 8610 24108
rect 8670 24108 8680 24120
rect 8582 24068 8594 24102
rect 8670 24068 8682 24108
rect 8582 24062 8682 24068
rect 8504 24040 8550 24052
rect 8504 23964 8510 24040
rect 8544 23964 8550 24040
rect 8714 24040 8760 24052
rect 8490 22964 8500 23964
rect 8552 23786 8562 23964
rect 8714 23963 8720 24040
rect 8754 23963 8760 24040
rect 8702 23786 8712 23963
rect 8552 22964 8712 23786
rect 8504 20072 8510 22964
rect 8544 22963 8712 22964
rect 8764 22963 8774 23963
rect 8544 20340 8720 22963
rect 8544 20072 8550 20340
rect 8504 20060 8550 20072
rect 8714 20072 8720 20340
rect 8754 20072 8760 22963
rect 8714 20060 8760 20072
rect 8582 20044 8682 20050
rect 8582 20004 8594 20044
rect 8670 20010 8682 20044
rect 8584 19992 8594 20004
rect 8654 20004 8682 20010
rect 8654 19992 8664 20004
rect 8852 19960 8858 24192
rect 8406 19954 8858 19960
rect 8892 24192 9344 24198
rect 8892 19960 8898 24192
rect 9070 24108 9080 24120
rect 9068 24068 9080 24108
rect 9140 24108 9150 24120
rect 9140 24102 9168 24108
rect 9156 24068 9168 24102
rect 9068 24062 9168 24068
rect 8990 24040 9036 24052
rect 8990 23963 8996 24040
rect 9030 23963 9036 24040
rect 9200 24040 9246 24052
rect 9200 23963 9206 24040
rect 9240 23963 9246 24040
rect 8977 22963 8987 23963
rect 9039 23786 9049 23963
rect 9187 23786 9197 23963
rect 9039 22963 9197 23786
rect 9249 22963 9259 23963
rect 8990 20072 8996 22963
rect 9030 20340 9206 22963
rect 9030 20072 9036 20340
rect 8990 20060 9036 20072
rect 9200 20072 9206 20340
rect 9240 20072 9246 22963
rect 9200 20060 9246 20072
rect 9068 20044 9168 20050
rect 9068 20010 9080 20044
rect 9068 20004 9096 20010
rect 9086 19992 9096 20004
rect 9156 20004 9168 20044
rect 9156 19992 9166 20004
rect 9338 19960 9344 24192
rect 8892 19954 9344 19960
rect 9378 24192 9830 24198
rect 9378 19960 9384 24192
rect 9572 24108 9582 24120
rect 9554 24102 9582 24108
rect 9642 24108 9652 24120
rect 9554 24068 9566 24102
rect 9642 24068 9654 24108
rect 9554 24062 9654 24068
rect 9476 24040 9522 24052
rect 9476 23963 9482 24040
rect 9516 23963 9522 24040
rect 9686 24040 9732 24052
rect 9686 23963 9692 24040
rect 9726 23963 9732 24040
rect 9463 22963 9473 23963
rect 9525 23786 9535 23963
rect 9674 23786 9684 23963
rect 9525 22963 9684 23786
rect 9736 22963 9746 23963
rect 9476 20072 9482 22963
rect 9516 20340 9692 22963
rect 9516 20072 9522 20340
rect 9476 20060 9522 20072
rect 9686 20072 9692 20340
rect 9726 20072 9732 22963
rect 9686 20060 9732 20072
rect 9554 20044 9654 20050
rect 9554 20004 9566 20044
rect 9642 20010 9654 20044
rect 9556 19992 9566 20004
rect 9626 20004 9654 20010
rect 9626 19992 9636 20004
rect 9824 19960 9830 24192
rect 9378 19954 9830 19960
rect 9864 24192 10316 24198
rect 9864 19960 9870 24192
rect 10042 24108 10052 24120
rect 10040 24068 10052 24108
rect 10112 24108 10122 24120
rect 10112 24102 10140 24108
rect 10128 24068 10140 24102
rect 10040 24062 10140 24068
rect 9962 24040 10008 24052
rect 9962 23963 9968 24040
rect 10002 23963 10008 24040
rect 10172 24040 10218 24052
rect 10172 23963 10178 24040
rect 10212 23963 10218 24040
rect 9949 22963 9959 23963
rect 10011 23786 10021 23963
rect 10159 23786 10169 23963
rect 10011 22963 10169 23786
rect 10221 22963 10231 23963
rect 9962 20072 9968 22963
rect 10002 20340 10178 22963
rect 10002 20072 10008 20340
rect 9962 20060 10008 20072
rect 10172 20072 10178 20340
rect 10212 20072 10218 22963
rect 10172 20060 10218 20072
rect 10040 20044 10140 20050
rect 10040 20010 10052 20044
rect 10040 20004 10068 20010
rect 10058 19992 10068 20004
rect 10128 20004 10140 20044
rect 10128 19992 10138 20004
rect 10310 19960 10316 24192
rect 9864 19954 10316 19960
rect 10350 24192 10771 24198
rect 10350 19960 10356 24192
rect 10544 24108 10554 24120
rect 10526 24102 10554 24108
rect 10614 24108 10624 24120
rect 10526 24068 10538 24102
rect 10614 24068 10626 24108
rect 10526 24062 10626 24068
rect 10448 24040 10494 24052
rect 10448 23963 10454 24040
rect 10488 23963 10494 24040
rect 10658 24040 10704 24052
rect 10436 22963 10446 23963
rect 10498 23789 10508 23963
rect 10658 23789 10664 24040
rect 10498 22963 10664 23789
rect 10448 20072 10454 22963
rect 10488 20343 10664 22963
rect 10488 20072 10494 20343
rect 10448 20060 10494 20072
rect 10658 20072 10664 20343
rect 10698 20072 10704 24040
rect 10658 20060 10704 20072
rect 10526 20044 10626 20050
rect 10526 20004 10538 20044
rect 10614 20010 10626 20044
rect 10528 19992 10538 20004
rect 10598 20004 10626 20010
rect 10598 19992 10608 20004
rect 10765 19960 10771 24192
rect 10855 24192 11244 24198
rect 10855 24189 10871 24192
rect 10855 23522 10861 24189
rect 15549 23843 15561 24198
rect 17598 24055 17610 24387
rect 19959 24055 20155 24061
rect 17598 24049 20155 24055
rect 15549 23837 15564 23843
rect 15552 23789 15564 23837
rect 15552 23783 19965 23789
rect 15847 23691 19839 23697
rect 15847 23657 15859 23691
rect 19827 23657 19839 23691
rect 15847 23651 19839 23657
rect 15791 23607 15837 23619
rect 10855 23516 10946 23522
rect 10855 23510 15607 23516
rect 15595 23364 15607 23510
rect 15778 23407 15788 23607
rect 15840 23407 15850 23607
rect 10918 23363 11074 23364
rect 10855 23358 11074 23363
rect 10855 23352 10946 23358
rect 10855 23351 10924 23352
rect 10855 20796 10861 23351
rect 11068 22337 11074 23358
rect 11220 23358 15607 23364
rect 11220 22362 11226 23358
rect 11341 23291 15383 23297
rect 11341 23257 11403 23291
rect 15371 23257 15383 23291
rect 11341 23251 15383 23257
rect 11341 23219 11375 23251
rect 11335 23207 11381 23219
rect 11335 22831 11341 23207
rect 11375 22831 11381 23207
rect 11322 22631 11332 22831
rect 11384 22631 11394 22831
rect 11335 22619 11381 22631
rect 11341 22587 11375 22619
rect 13036 22587 13886 23251
rect 15393 23207 15439 23219
rect 15393 22831 15399 23207
rect 15433 22831 15439 23207
rect 15380 22631 15390 22831
rect 15442 22631 15452 22831
rect 15791 22631 15797 23407
rect 15831 22631 15837 23407
rect 15393 22619 15439 22631
rect 15791 22619 15837 22631
rect 17472 22587 18326 23651
rect 19849 23607 19895 23619
rect 19836 23407 19846 23607
rect 19898 23407 19908 23607
rect 19849 22631 19855 23407
rect 19889 22631 19895 23407
rect 19849 22619 19895 22631
rect 11341 22581 19839 22587
rect 11341 22547 11403 22581
rect 15371 22547 15859 22581
rect 19827 22547 19839 22581
rect 11341 22541 19839 22547
rect 15183 22478 16047 22541
rect 11220 22356 15138 22362
rect 11068 22172 11080 22337
rect 15126 22172 15138 22356
rect 11068 22166 11200 22172
rect 10855 20790 10869 20796
rect 11194 20790 11200 22166
rect 10855 20784 11200 20790
rect 11261 22166 15138 22172
rect 11261 20790 11267 22166
rect 15183 22088 15383 22478
rect 15847 22088 16047 22478
rect 19959 22393 19965 23783
rect 16135 22387 19965 22393
rect 16135 22146 16147 22387
rect 16135 22140 19965 22146
rect 15183 22025 16047 22088
rect 11398 22019 19839 22025
rect 11398 21985 11410 22019
rect 15378 21985 15859 22019
rect 19827 21985 19839 22019
rect 11398 21979 19839 21985
rect 11342 21935 11388 21947
rect 11342 21159 11348 21935
rect 11382 21159 11388 21935
rect 11329 20959 11339 21159
rect 11391 20959 11401 21159
rect 11342 20947 11388 20959
rect 13025 20915 13879 21979
rect 15797 21947 15831 21979
rect 15400 21935 15446 21947
rect 15791 21935 15837 21947
rect 15400 21159 15406 21935
rect 15440 21159 15446 21935
rect 15524 21768 15692 21780
rect 15520 21161 15530 21768
rect 15686 21195 15696 21768
rect 15778 21735 15788 21935
rect 15840 21735 15850 21935
rect 15791 21359 15797 21735
rect 15831 21359 15837 21735
rect 15791 21347 15837 21359
rect 15797 21315 15831 21347
rect 17497 21315 18347 21979
rect 19849 21935 19895 21947
rect 19836 21735 19846 21935
rect 19898 21735 19908 21935
rect 19959 21752 19965 22140
rect 20149 21752 20155 24049
rect 19849 21359 19855 21735
rect 19889 21359 19895 21735
rect 19849 21347 19895 21359
rect 15797 21309 19839 21315
rect 15797 21275 15859 21309
rect 19827 21275 19839 21309
rect 15797 21269 19839 21275
rect 19951 21195 19961 21752
rect 15686 21189 19961 21195
rect 15387 20959 15397 21159
rect 15449 20959 15459 21159
rect 15520 21075 15532 21161
rect 20149 21110 20158 21752
rect 20149 21081 20155 21110
rect 15400 20947 15446 20959
rect 11398 20909 15390 20915
rect 11398 20875 11410 20909
rect 15378 20875 15390 20909
rect 11398 20869 15390 20875
rect 11261 20789 11275 20790
rect 15526 20789 15532 21075
rect 11261 20784 15532 20789
rect 11263 20783 15532 20784
rect 15600 21075 20155 21081
rect 15600 20789 15606 21075
rect 19959 21069 20155 21075
rect 15600 20783 15615 20789
rect 15603 20696 15615 20783
rect 10350 19954 10771 19960
rect 10855 20690 15615 20696
rect 10855 20684 10869 20690
rect 11194 20684 11267 20690
rect 15526 20687 15606 20690
rect 10855 19739 10861 20684
rect 10825 19731 10861 19739
rect 5730 19727 10861 19731
rect 5730 19725 10837 19727
rect 6135 19372 6258 19378
rect 19965 19372 20101 19378
rect 6135 19366 20106 19372
rect 6135 16881 6141 19366
rect 6124 16875 6141 16881
rect 6252 19240 10574 19246
rect 6252 16881 6258 19240
rect 9340 19138 9350 19143
rect 6408 19132 9350 19138
rect 10350 19138 10360 19143
rect 10350 19132 10404 19138
rect 6408 19098 6420 19132
rect 10388 19098 10404 19132
rect 6408 19092 9350 19098
rect 6743 19087 9350 19092
rect 10350 19092 10404 19098
rect 10350 19087 10360 19092
rect 6352 19039 6398 19051
rect 6339 18763 6349 19039
rect 6401 18763 6411 19039
rect 6352 18751 6398 18763
rect 6743 18710 10119 19087
rect 10410 19039 10456 19051
rect 10397 18763 10407 19039
rect 10459 18763 10469 19039
rect 10410 18751 10456 18763
rect 6408 18704 10400 18710
rect 6408 18670 6420 18704
rect 10388 18670 10400 18704
rect 6408 18664 10400 18670
rect 6514 18602 10365 18664
rect 6408 18596 10400 18602
rect 6408 18562 6420 18596
rect 10388 18562 10400 18596
rect 6408 18556 10400 18562
rect 6352 18503 6398 18515
rect 6339 18227 6349 18503
rect 6401 18227 6411 18503
rect 6352 18215 6398 18227
rect 6738 18174 10108 18556
rect 10410 18503 10456 18515
rect 10397 18227 10407 18503
rect 10459 18227 10469 18503
rect 10410 18215 10456 18227
rect 6408 18168 10400 18174
rect 6408 18134 6420 18168
rect 10388 18134 10400 18168
rect 6408 18128 10400 18134
rect 9912 17738 10291 18128
rect 6408 17732 10400 17738
rect 6408 17698 6420 17732
rect 10388 17698 10400 17732
rect 6408 17692 10400 17698
rect 6352 17639 6398 17651
rect 6332 17439 6342 17639
rect 6406 17439 6416 17639
rect 6352 17063 6358 17439
rect 6392 17063 6398 17439
rect 6352 17051 6398 17063
rect 6666 17010 10039 17692
rect 10410 17639 10456 17651
rect 10397 17063 10407 17639
rect 10459 17063 10469 17639
rect 10410 17051 10456 17063
rect 6408 17004 10404 17010
rect 6408 16970 6420 17004
rect 10388 16970 10404 17004
rect 6408 16964 10404 16970
rect 7981 16881 8249 16886
rect 10568 16881 10574 19240
rect 6252 16875 10574 16881
rect 11339 19240 19971 19246
rect 6124 16741 6136 16875
rect 6124 16735 8056 16741
rect 6135 16733 6258 16735
rect 8050 14789 8056 16735
rect 8243 15035 10574 15041
rect 8243 14789 8249 15035
rect 8410 14885 8420 14937
rect 9420 14934 9430 14937
rect 9420 14928 10400 14934
rect 10388 14894 10400 14928
rect 9420 14888 10400 14894
rect 9420 14885 10204 14888
rect 8362 14835 8408 14847
rect 8044 14450 8054 14789
rect 8246 14470 8256 14789
rect 8362 14786 8368 14835
rect 8402 14786 8408 14835
rect 8339 14659 8349 14786
rect 8402 14659 8411 14786
rect 8362 14647 8408 14659
rect 8683 14606 10204 14885
rect 10410 14835 10456 14847
rect 10397 14659 10407 14835
rect 10459 14659 10469 14835
rect 10410 14647 10456 14659
rect 8418 14600 10400 14606
rect 8418 14566 8430 14600
rect 10388 14566 10400 14600
rect 8418 14560 10400 14566
rect 10568 14470 10574 15035
rect 8246 14464 10574 14470
rect 11339 14470 11345 19240
rect 11496 19138 11506 19143
rect 11492 19092 11506 19138
rect 12506 19138 12516 19143
rect 12506 19132 19870 19138
rect 15476 19098 15834 19132
rect 19802 19098 19870 19132
rect 11496 19087 11506 19092
rect 12506 19092 19870 19098
rect 12506 19087 12516 19092
rect 11440 19039 11486 19051
rect 11440 17663 11446 19039
rect 11480 17663 11486 19039
rect 11421 17063 11431 17663
rect 11495 17063 11505 17663
rect 11440 17051 11486 17063
rect 13053 17010 14232 19092
rect 15498 19039 15544 19051
rect 15498 17563 15504 19039
rect 15538 18929 15544 19039
rect 15766 19039 15812 19051
rect 15766 18929 15772 19039
rect 15538 17563 15772 18929
rect 15806 17563 15812 19039
rect 15485 17063 15495 17563
rect 15547 17155 15763 17563
rect 15547 17063 15557 17155
rect 15753 17063 15763 17155
rect 15815 17063 15825 17563
rect 15498 17051 15544 17063
rect 15766 17051 15812 17063
rect 17305 17010 18484 19092
rect 19824 19039 19870 19092
rect 19805 18439 19815 19039
rect 19879 18439 19889 19039
rect 19965 18903 19971 19240
rect 20095 19240 20106 19366
rect 20095 18995 20101 19240
rect 20564 18995 21843 18998
rect 20095 18992 21843 18995
rect 20095 18983 20576 18992
rect 19965 18891 19989 18903
rect 19824 17063 19830 18439
rect 19864 17063 19870 18439
rect 19824 17051 19870 17063
rect 19830 17010 19864 17051
rect 11492 17004 19864 17010
rect 11492 16970 11508 17004
rect 15476 16970 15834 17004
rect 19802 16970 19864 17004
rect 11492 16964 19864 16970
rect 11505 16734 15414 16964
rect 15894 16734 19803 16964
rect 11440 16728 19814 16734
rect 11440 16694 11508 16728
rect 15476 16694 15834 16728
rect 19802 16694 19814 16728
rect 11440 16688 19814 16694
rect 11440 16635 11486 16688
rect 11421 16035 11431 16635
rect 11495 16035 11505 16635
rect 11440 14659 11446 16035
rect 11480 14659 11486 16035
rect 11440 14647 11486 14659
rect 11446 14606 11486 14647
rect 13019 14606 14198 16688
rect 15498 16635 15544 16647
rect 15766 16635 15812 16647
rect 15485 16135 15495 16635
rect 15547 16531 15557 16635
rect 15753 16531 15763 16635
rect 15547 16135 15763 16531
rect 15815 16135 15825 16635
rect 15498 14850 15504 16135
rect 15538 14850 15772 16135
rect 15806 14850 15812 16135
rect 15485 14659 15495 14850
rect 15547 14745 15763 14850
rect 15547 14659 15557 14745
rect 15753 14659 15763 14745
rect 15815 14659 15825 14850
rect 15498 14647 15544 14659
rect 15766 14647 15812 14659
rect 17322 14606 18501 16688
rect 19824 16635 19870 16647
rect 19824 15259 19830 16635
rect 19864 15259 19870 16635
rect 19805 14792 19815 15259
rect 19879 14792 19889 15259
rect 19805 14778 19830 14792
rect 19824 14659 19830 14778
rect 19864 14778 19889 14792
rect 19864 14659 19870 14778
rect 19824 14647 19870 14659
rect 11446 14600 19814 14606
rect 11446 14566 11508 14600
rect 15476 14566 15834 14600
rect 19802 14566 19814 14600
rect 11446 14560 19814 14566
rect 19983 14470 19989 18891
rect 21831 18859 21843 18992
rect 11339 14464 19989 14470
rect 20718 18853 21688 18859
rect 20718 14470 20724 18853
rect 20901 18774 20911 18780
rect 20899 18728 20911 18774
rect 20987 18774 20997 18780
rect 20987 18728 20999 18774
rect 21393 18732 21403 18796
rect 21503 18732 21513 18796
rect 21403 18728 21503 18732
rect 20812 18706 20858 18718
rect 20812 14738 20818 18706
rect 20852 18069 20858 18706
rect 21040 18706 21086 18718
rect 21040 18700 21046 18706
rect 21080 18700 21086 18706
rect 21316 18706 21362 18718
rect 21025 18069 21035 18700
rect 20852 17700 21035 18069
rect 21091 17700 21101 18700
rect 20852 15472 21046 17700
rect 20852 14738 20858 15472
rect 20812 14726 20858 14738
rect 21040 14738 21046 15472
rect 21080 14738 21086 17700
rect 21040 14726 21086 14738
rect 21316 14738 21322 18706
rect 21356 18069 21362 18706
rect 21544 18706 21590 18718
rect 21544 18658 21550 18706
rect 21584 18658 21590 18706
rect 21529 18069 21539 18658
rect 21356 17658 21539 18069
rect 21595 17658 21605 18658
rect 21356 15472 21550 17658
rect 21356 14738 21362 15472
rect 21316 14726 21362 14738
rect 21544 14738 21550 15472
rect 21584 14738 21590 17658
rect 21544 14726 21590 14738
rect 20899 14670 20911 14716
rect 20901 14664 20911 14670
rect 20987 14670 20999 14716
rect 21403 14670 21415 14716
rect 20987 14664 20997 14670
rect 21405 14664 21415 14670
rect 21491 14670 21503 14716
rect 21491 14664 21501 14670
rect 21682 14470 21688 18853
rect 20718 14464 21688 14470
rect 21822 18853 21843 18859
rect 21822 14454 21828 18853
rect 8044 14001 8056 14450
rect 8044 13995 21564 14001
rect 21554 13991 21564 13995
rect 21822 13991 21832 14454
rect 7788 12824 10790 12830
rect 7788 12572 7800 12824
rect 10778 12663 10790 12824
rect 7788 12513 7796 12572
rect 5834 11975 5989 11981
rect 7790 11975 7796 12513
rect 5834 11969 7796 11975
rect 7999 12513 10284 12519
rect 7999 11975 8005 12513
rect 8123 12404 10125 12410
rect 8123 12370 8135 12404
rect 10113 12370 10125 12404
rect 8123 12364 10125 12370
rect 8054 12135 8064 12335
rect 8116 12135 8126 12335
rect 8067 12123 8113 12135
rect 8436 12084 9785 12364
rect 10135 12311 10181 12323
rect 10112 12135 10122 12311
rect 10175 12135 10184 12311
rect 10135 12123 10181 12135
rect 8125 12082 8135 12084
rect 8123 12036 8135 12082
rect 8844 12082 9785 12084
rect 8844 12076 10125 12082
rect 10113 12042 10125 12076
rect 8125 12032 8135 12036
rect 8844 12036 10125 12042
rect 8844 12032 8854 12036
rect 10274 11975 10284 12513
rect 7999 11969 10284 11975
rect 5826 11194 5836 11969
rect 5983 11751 10284 11757
rect 5983 11194 5993 11751
rect 6123 11641 10115 11647
rect 6123 11607 6135 11641
rect 10103 11607 10115 11641
rect 6123 11601 10115 11607
rect 6067 11548 6113 11560
rect 5834 10956 5840 11194
rect 5983 10988 5989 11194
rect 6048 11172 6058 11548
rect 6116 11172 6126 11548
rect 6067 11160 6113 11172
rect 7025 11119 9474 11601
rect 10125 11548 10171 11560
rect 10112 11172 10122 11548
rect 10174 11172 10184 11548
rect 10125 11160 10171 11172
rect 6123 11115 10115 11119
rect 6123 11073 6135 11115
rect 7135 11113 10115 11115
rect 10103 11079 10115 11113
rect 6125 11063 6135 11073
rect 7135 11073 10115 11079
rect 7135 11063 7145 11073
rect 10274 10988 10284 11751
rect 5983 10982 10284 10988
rect 5830 10840 5840 10956
rect 5834 10801 5840 10840
rect 5834 10789 5844 10801
rect 5838 8767 5844 10789
rect 6065 10795 7787 10801
rect 6065 8877 6071 10795
rect 6235 10655 6707 10661
rect 6235 10621 6247 10655
rect 6695 10621 6707 10655
rect 6235 10615 6707 10621
rect 7171 10655 7643 10661
rect 7171 10621 7183 10655
rect 7631 10621 7643 10655
rect 7171 10615 7643 10621
rect 6179 10562 6225 10574
rect 6160 10327 6170 10562
rect 6234 10327 6244 10562
rect 6179 10086 6185 10327
rect 6219 10086 6225 10327
rect 6179 10074 6225 10086
rect 6366 10033 6558 10615
rect 6717 10562 6763 10574
rect 6717 10086 6723 10562
rect 6757 10192 6763 10562
rect 7115 10562 7161 10574
rect 6882 10192 6892 10194
rect 6757 10086 6892 10192
rect 6717 10074 6892 10086
rect 6235 10027 6707 10033
rect 6235 9993 6247 10027
rect 6695 9993 6707 10027
rect 6235 9987 6707 9993
rect 6235 9918 6335 9987
rect 6882 9970 6892 10074
rect 6985 10192 6995 10194
rect 7115 10192 7121 10562
rect 6985 10086 7121 10192
rect 7155 10086 7161 10562
rect 6985 10074 7161 10086
rect 6985 9970 6995 10074
rect 7313 10033 7505 10615
rect 7653 10562 7699 10574
rect 7653 10322 7659 10562
rect 7693 10322 7699 10562
rect 7634 10086 7644 10322
rect 7708 10086 7718 10322
rect 7653 10074 7699 10086
rect 7171 10027 7643 10033
rect 7171 9993 7183 10027
rect 7631 9993 7643 10027
rect 7171 9987 7649 9993
rect 6225 9818 6235 9918
rect 6335 9818 6345 9918
rect 6597 9668 6607 9768
rect 6707 9668 6717 9768
rect 6607 9619 6707 9668
rect 6235 9613 6707 9619
rect 6235 9579 6247 9613
rect 6695 9579 6707 9613
rect 6235 9573 6707 9579
rect 6179 9520 6225 9532
rect 6179 9280 6185 9520
rect 6219 9280 6225 9520
rect 6160 9044 6170 9280
rect 6234 9044 6244 9280
rect 6179 9032 6225 9044
rect 6366 8991 6558 9573
rect 6886 9532 6986 9970
rect 7161 9818 7171 9918
rect 7271 9818 7281 9918
rect 7171 9619 7271 9818
rect 7549 9768 7649 9987
rect 7539 9668 7549 9768
rect 7649 9668 7659 9768
rect 7171 9613 7643 9619
rect 7171 9579 7183 9613
rect 7631 9579 7643 9613
rect 7171 9573 7643 9579
rect 6717 9520 7161 9532
rect 6717 9044 6723 9520
rect 6757 9414 7121 9520
rect 6757 9044 6763 9414
rect 6717 9032 6763 9044
rect 7115 9044 7121 9414
rect 7155 9044 7161 9520
rect 7115 9032 7161 9044
rect 7308 8991 7500 9573
rect 7653 9520 7699 9532
rect 7634 9285 7644 9520
rect 7708 9285 7718 9520
rect 7653 9044 7659 9285
rect 7693 9044 7699 9285
rect 7653 9032 7699 9044
rect 6235 8985 6707 8991
rect 6235 8951 6247 8985
rect 6695 8951 6707 8985
rect 6235 8945 6707 8951
rect 7171 8985 7643 8991
rect 7171 8951 7183 8985
rect 7631 8951 7643 8985
rect 7171 8945 7643 8951
rect 7777 8877 7787 10795
rect 6065 8871 7787 8877
rect 7942 10795 8812 10801
rect 7942 8877 7952 10795
rect 7942 8871 7972 8877
rect 7960 8767 7972 8871
rect 5838 8761 7972 8767
rect 5838 8755 6071 8761
rect 8802 8741 8812 10795
rect 10779 12513 10790 12663
rect 10779 10806 10789 12513
rect 11842 11123 11973 11126
rect 11842 11117 12911 11123
rect 11842 11114 11880 11117
rect 10361 10801 10655 10806
rect 8950 10795 10655 10801
rect 8950 8869 8960 10795
rect 10278 10794 10655 10795
rect 9101 10673 9573 10679
rect 9101 10639 9113 10673
rect 9561 10639 9573 10673
rect 9101 10633 9573 10639
rect 10033 10673 10555 10679
rect 10033 10639 10045 10673
rect 10493 10639 10555 10673
rect 10033 10633 10555 10639
rect 9045 10580 9091 10592
rect 9045 10304 9051 10580
rect 9085 10304 9091 10580
rect 9026 10104 9036 10304
rect 9100 10104 9110 10304
rect 9045 10092 9091 10104
rect 9193 10051 9444 10633
rect 9583 10580 9629 10592
rect 9977 10580 10023 10592
rect 9570 10380 9580 10580
rect 9632 10380 9642 10580
rect 9964 10380 9974 10580
rect 10026 10380 10036 10580
rect 9583 10104 9589 10380
rect 9623 10104 9629 10380
rect 9583 10092 9629 10104
rect 9977 10104 9983 10380
rect 10017 10104 10023 10380
rect 9977 10092 10023 10104
rect 10166 10051 10374 10633
rect 10521 10592 10555 10633
rect 10515 10580 10561 10592
rect 10496 10380 10506 10580
rect 10570 10380 10580 10580
rect 10515 10104 10521 10380
rect 10555 10104 10561 10380
rect 10515 10092 10561 10104
rect 10521 10051 10555 10092
rect 9101 10045 9573 10051
rect 10033 10045 10555 10051
rect 9101 10011 9113 10045
rect 9561 10011 10045 10045
rect 10493 10011 10555 10045
rect 9101 10005 9573 10011
rect 9448 9594 9573 10005
rect 9051 9588 9573 9594
rect 10033 10005 10555 10011
rect 10033 9594 10158 10005
rect 10033 9588 10505 9594
rect 9051 9554 9113 9588
rect 9561 9554 10045 9588
rect 10493 9554 10505 9588
rect 9051 9548 9573 9554
rect 10033 9548 10505 9554
rect 9051 9507 9085 9548
rect 9045 9495 9091 9507
rect 9026 9295 9036 9495
rect 9100 9295 9110 9495
rect 9045 9019 9051 9295
rect 9085 9019 9091 9295
rect 9045 9007 9091 9019
rect 9051 8966 9085 9007
rect 9236 8966 9444 9548
rect 9583 9495 9629 9507
rect 9977 9495 10023 9507
rect 9570 9295 9580 9495
rect 9632 9295 9642 9495
rect 9964 9295 9974 9495
rect 10026 9295 10036 9495
rect 9583 9019 9589 9295
rect 9623 9019 9629 9295
rect 9583 9007 9629 9019
rect 9977 9019 9983 9295
rect 10017 9019 10023 9295
rect 9977 9007 10023 9019
rect 10153 8966 10361 9548
rect 10515 9495 10561 9507
rect 10515 9219 10521 9495
rect 10555 9219 10561 9495
rect 10496 9019 10506 9219
rect 10570 9019 10580 9219
rect 10515 9007 10561 9019
rect 9051 8960 9573 8966
rect 9051 8926 9113 8960
rect 9561 8926 9573 8960
rect 9051 8920 9573 8926
rect 10033 8960 10505 8966
rect 10033 8926 10045 8960
rect 10493 8926 10505 8960
rect 10033 8920 10505 8926
rect 10645 8869 10655 10794
rect 8950 8863 10655 8869
rect 8806 8737 8821 8741
rect 8806 8731 10655 8737
rect 8806 8729 8956 8731
rect 10645 8728 10655 8731
rect 10776 8728 10786 10806
rect 11838 10404 11848 11114
rect 12899 11079 12911 11117
rect 11967 11000 12773 11006
rect 11967 10404 11977 11000
rect 12083 10946 12175 10952
rect 12083 10912 12095 10946
rect 12163 10912 12175 10946
rect 12083 10906 12175 10912
rect 12241 10946 12333 10952
rect 12241 10912 12253 10946
rect 12321 10912 12333 10946
rect 12241 10906 12333 10912
rect 12399 10946 12491 10952
rect 12399 10912 12411 10946
rect 12479 10912 12491 10946
rect 12399 10906 12491 10912
rect 12557 10946 12649 10952
rect 12557 10912 12569 10946
rect 12637 10912 12649 10946
rect 12557 10906 12649 10912
rect 12027 10853 12073 10865
rect 12027 10777 12033 10853
rect 12067 10777 12073 10853
rect 12014 10677 12024 10777
rect 12076 10677 12086 10777
rect 12027 10665 12073 10677
rect 12115 10624 12151 10906
rect 12265 10905 12301 10906
rect 12185 10853 12231 10865
rect 12185 10677 12191 10853
rect 12225 10677 12231 10853
rect 12185 10665 12231 10677
rect 12266 10625 12299 10905
rect 12343 10853 12389 10865
rect 12330 10753 12340 10853
rect 12392 10753 12402 10853
rect 12343 10677 12349 10753
rect 12383 10677 12389 10753
rect 12343 10665 12389 10677
rect 12265 10624 12301 10625
rect 12430 10624 12466 10906
rect 12501 10853 12547 10865
rect 12501 10677 12507 10853
rect 12541 10677 12547 10853
rect 12501 10665 12547 10677
rect 12582 10624 12618 10906
rect 12659 10853 12705 10865
rect 12659 10777 12665 10853
rect 12699 10777 12705 10853
rect 12646 10677 12656 10777
rect 12708 10677 12718 10777
rect 12659 10665 12705 10677
rect 12083 10618 12175 10624
rect 12083 10584 12095 10618
rect 12163 10584 12175 10618
rect 12083 10578 12175 10584
rect 12241 10618 12333 10624
rect 12241 10584 12253 10618
rect 12321 10584 12333 10618
rect 12241 10578 12333 10584
rect 12399 10618 12491 10624
rect 12399 10584 12411 10618
rect 12479 10584 12491 10618
rect 12399 10578 12491 10584
rect 12557 10618 12649 10624
rect 12557 10584 12569 10618
rect 12637 10584 12649 10618
rect 12557 10578 12649 10584
rect 11842 10392 11973 10404
rect 12083 10349 12133 10578
rect 12083 10295 12148 10349
rect 12203 10295 12213 10349
rect 12083 10113 12133 10295
rect 11509 10063 12133 10113
rect 11235 9898 11316 9910
rect 11231 9293 11241 9898
rect 11229 9173 11241 9293
rect 11310 9293 11320 9898
rect 11509 9728 11559 10063
rect 12241 10015 12291 10578
rect 12399 10226 12449 10578
rect 12320 10172 12330 10226
rect 12384 10172 12449 10226
rect 12065 9965 12291 10015
rect 12399 10015 12449 10172
rect 12557 10113 12607 10578
rect 12763 10418 12773 11000
rect 12901 10418 12911 11079
rect 13747 11048 13879 11054
rect 13747 11042 20429 11048
rect 13747 11032 13753 11042
rect 12767 10406 12907 10418
rect 12557 10063 13185 10113
rect 12399 9965 12629 10015
rect 11467 9722 11559 9728
rect 11467 9688 11479 9722
rect 11547 9688 11559 9722
rect 11467 9682 11559 9688
rect 11717 9898 11854 9910
rect 11411 9638 11457 9650
rect 11569 9638 11615 9650
rect 11398 9558 11408 9638
rect 11460 9558 11470 9638
rect 11411 9462 11417 9558
rect 11451 9462 11457 9558
rect 11569 9542 11575 9638
rect 11609 9542 11615 9638
rect 11556 9462 11566 9542
rect 11618 9462 11628 9542
rect 11411 9450 11457 9462
rect 11569 9450 11615 9462
rect 11467 9412 11559 9418
rect 11467 9378 11479 9412
rect 11547 9378 11559 9412
rect 11467 9372 11559 9378
rect 11717 9293 11723 9898
rect 11310 9287 11723 9293
rect 11848 9293 11854 9898
rect 12065 9728 12115 9965
rect 12023 9722 12115 9728
rect 12023 9688 12035 9722
rect 12103 9688 12115 9722
rect 12023 9682 12115 9688
rect 12274 9901 12411 9913
rect 11967 9638 12013 9650
rect 12125 9638 12171 9650
rect 11967 9542 11973 9638
rect 12007 9542 12013 9638
rect 12112 9558 12122 9638
rect 12174 9558 12184 9638
rect 11954 9462 11964 9542
rect 12016 9462 12026 9542
rect 12125 9462 12131 9558
rect 12165 9462 12171 9558
rect 11967 9450 12013 9462
rect 12125 9450 12171 9462
rect 12023 9412 12115 9418
rect 12023 9372 12035 9412
rect 12025 9356 12035 9372
rect 12103 9372 12115 9412
rect 12103 9356 12113 9372
rect 12274 9293 12280 9901
rect 11848 9287 12280 9293
rect 12405 9293 12411 9901
rect 12579 9728 12629 9965
rect 12838 9893 12975 9905
rect 12579 9722 12671 9728
rect 12579 9688 12591 9722
rect 12659 9688 12671 9722
rect 12579 9682 12671 9688
rect 12523 9638 12569 9650
rect 12681 9638 12727 9650
rect 12510 9558 12520 9638
rect 12572 9558 12582 9638
rect 12523 9462 12529 9558
rect 12563 9462 12569 9558
rect 12681 9542 12687 9638
rect 12721 9542 12727 9638
rect 12668 9462 12678 9542
rect 12730 9462 12740 9542
rect 12523 9450 12569 9462
rect 12681 9450 12727 9462
rect 12579 9412 12671 9418
rect 12579 9378 12591 9412
rect 12659 9378 12671 9412
rect 12579 9372 12671 9378
rect 12838 9293 12844 9893
rect 12405 9287 12844 9293
rect 12969 9293 12975 9893
rect 13135 9728 13185 10063
rect 13378 9900 13454 9912
rect 13135 9722 13227 9728
rect 13135 9688 13147 9722
rect 13215 9688 13227 9722
rect 13135 9682 13227 9688
rect 13079 9638 13125 9650
rect 13237 9638 13283 9650
rect 13079 9542 13085 9638
rect 13119 9542 13125 9638
rect 13224 9558 13234 9638
rect 13286 9558 13296 9638
rect 13066 9462 13076 9542
rect 13128 9462 13138 9542
rect 13237 9462 13243 9558
rect 13277 9462 13283 9558
rect 13079 9450 13125 9462
rect 13237 9450 13283 9462
rect 13135 9412 13227 9418
rect 13135 9372 13147 9412
rect 13137 9356 13147 9372
rect 13215 9372 13227 9412
rect 13215 9356 13225 9372
rect 13374 9293 13384 9900
rect 12969 9287 13384 9293
rect 13448 9287 13458 9900
rect 13446 9173 13458 9287
rect 11229 9167 13458 9173
rect 10649 8716 10782 8728
rect 8517 8650 8595 8662
rect 8513 8646 8523 8650
rect 5306 8642 8523 8646
rect 5289 8640 8523 8642
rect 5289 8630 5318 8640
rect 8589 8632 8599 8650
rect 5285 5730 5295 8630
rect 8589 8626 10802 8632
rect 5375 8554 8523 8560
rect 5375 8015 5385 8554
rect 5515 8471 6707 8477
rect 7171 8471 8363 8477
rect 5465 8437 5527 8471
rect 6695 8437 7183 8471
rect 8351 8437 8363 8471
rect 5465 8431 6707 8437
rect 7171 8431 8363 8437
rect 5465 8399 5499 8431
rect 5459 8387 5505 8399
rect 6717 8387 6763 8399
rect 7115 8387 7161 8399
rect 8373 8387 8419 8399
rect 5440 8323 5450 8387
rect 5514 8323 5524 8387
rect 5459 8211 5465 8323
rect 5499 8211 5505 8323
rect 6704 8287 6714 8387
rect 6766 8287 6776 8387
rect 7102 8287 7112 8387
rect 7164 8287 7174 8387
rect 5459 8199 5505 8211
rect 6717 8211 6723 8287
rect 6757 8211 6763 8287
rect 6717 8199 6763 8211
rect 7115 8211 7121 8287
rect 7155 8211 7161 8287
rect 8373 8275 8379 8387
rect 8413 8275 8419 8387
rect 8354 8211 8364 8275
rect 8428 8211 8438 8275
rect 7115 8199 7161 8211
rect 8373 8199 8419 8211
rect 5464 8167 5499 8199
rect 5464 8161 6707 8167
rect 7171 8161 8363 8167
rect 5464 8127 5527 8161
rect 6695 8127 7183 8161
rect 8351 8127 8363 8161
rect 5464 8121 6707 8127
rect 7171 8121 8363 8127
rect 8513 8015 8523 8554
rect 5375 8009 8523 8015
rect 8589 8558 8824 8564
rect 8589 8001 8599 8558
rect 8814 8001 8824 8558
rect 8589 7995 8824 8001
rect 8961 8558 9704 8564
rect 8961 8001 8971 8558
rect 9101 8471 9533 8477
rect 9101 8437 9113 8471
rect 9521 8437 9533 8471
rect 9101 8431 9533 8437
rect 9045 8387 9091 8399
rect 9543 8387 9589 8399
rect 9026 8287 9036 8387
rect 9100 8287 9110 8387
rect 9543 8311 9549 8387
rect 9583 8311 9589 8387
rect 9045 8211 9051 8287
rect 9085 8211 9091 8287
rect 9530 8211 9540 8311
rect 9592 8211 9602 8311
rect 9045 8199 9091 8211
rect 9543 8199 9589 8211
rect 9103 8167 9113 8171
rect 9101 8121 9113 8167
rect 9273 8167 9283 8171
rect 9273 8161 9533 8167
rect 9521 8127 9533 8161
rect 9103 8107 9113 8121
rect 9273 8121 9533 8127
rect 9273 8107 9283 8121
rect 9694 8001 9704 8558
rect 8961 7995 9704 8001
rect 9897 8558 10665 8564
rect 9897 8001 9907 8558
rect 10073 8472 10505 8478
rect 10073 8438 10085 8472
rect 10493 8438 10505 8472
rect 10073 8432 10505 8438
rect 10017 8388 10063 8400
rect 10515 8388 10561 8400
rect 10004 8288 10014 8388
rect 10066 8288 10076 8388
rect 10496 8288 10506 8388
rect 10570 8288 10580 8388
rect 10017 8212 10023 8288
rect 10057 8212 10063 8288
rect 10017 8200 10063 8212
rect 10515 8212 10521 8288
rect 10555 8212 10561 8288
rect 10515 8200 10561 8212
rect 10075 8168 10085 8173
rect 10073 8122 10085 8168
rect 10245 8168 10255 8173
rect 10245 8162 10505 8168
rect 10493 8128 10505 8162
rect 10075 8109 10085 8122
rect 10245 8122 10505 8128
rect 10245 8109 10255 8122
rect 10655 8001 10665 8558
rect 9897 7995 10665 8001
rect 10790 8558 10802 8626
rect 10790 8001 10800 8558
rect 10790 7995 10814 8001
rect 10802 7933 10814 7995
rect 8589 7927 10814 7933
rect 5375 7863 8523 7869
rect 5375 7301 5385 7863
rect 5465 7755 6707 7761
rect 7171 7755 8363 7761
rect 5465 7721 5527 7755
rect 6695 7721 7183 7755
rect 8351 7721 8363 7755
rect 5465 7715 6707 7721
rect 7171 7715 8363 7721
rect 5465 7683 5499 7715
rect 5459 7671 5505 7683
rect 6717 7671 6763 7683
rect 5440 7607 5450 7671
rect 5514 7607 5524 7671
rect 5459 7495 5465 7607
rect 5499 7495 5505 7607
rect 6717 7595 6723 7671
rect 6757 7595 6763 7671
rect 7115 7671 7161 7683
rect 7115 7595 7121 7671
rect 7155 7595 7161 7671
rect 8373 7671 8419 7683
rect 6704 7495 6714 7595
rect 6766 7495 6776 7595
rect 7102 7495 7112 7595
rect 7164 7495 7174 7595
rect 8373 7548 8379 7671
rect 8413 7548 8419 7671
rect 5459 7483 5505 7495
rect 6717 7483 6763 7495
rect 7115 7483 7161 7495
rect 8354 7484 8364 7548
rect 8428 7484 8438 7548
rect 8373 7483 8419 7484
rect 5465 7451 5499 7483
rect 5465 7445 6707 7451
rect 7171 7445 8363 7451
rect 5465 7411 5527 7445
rect 6695 7411 7183 7445
rect 8351 7411 8363 7445
rect 5465 7405 6707 7411
rect 7171 7405 8363 7411
rect 8513 7301 8523 7863
rect 5375 7295 8523 7301
rect 5375 7149 8523 7155
rect 5375 6570 5385 7149
rect 5515 7039 6707 7045
rect 7171 7039 8413 7045
rect 5515 7005 5527 7039
rect 6695 7005 7183 7039
rect 8351 7005 8413 7039
rect 5515 6999 6707 7005
rect 7171 6999 8413 7005
rect 8379 6967 8413 6999
rect 5459 6955 5505 6967
rect 6717 6955 6763 6967
rect 5440 6891 5450 6955
rect 5514 6891 5524 6955
rect 5459 6779 5465 6891
rect 5499 6779 5505 6891
rect 6717 6879 6723 6955
rect 6757 6879 6763 6955
rect 7115 6955 7161 6967
rect 8373 6955 8419 6967
rect 7115 6879 7121 6955
rect 7155 6879 7161 6955
rect 8354 6891 8364 6955
rect 8428 6891 8438 6955
rect 6704 6779 6714 6879
rect 6766 6779 6776 6879
rect 7102 6779 7112 6879
rect 7164 6779 7174 6879
rect 8373 6779 8379 6891
rect 8413 6779 8419 6891
rect 5459 6767 5505 6779
rect 6717 6767 6763 6779
rect 7115 6767 7161 6779
rect 8373 6767 8419 6779
rect 8379 6735 8413 6767
rect 5515 6729 6707 6735
rect 7171 6729 8413 6735
rect 5515 6695 5527 6729
rect 6695 6695 7183 6729
rect 8351 6695 8413 6729
rect 5515 6689 6707 6695
rect 7171 6689 8413 6695
rect 8513 6570 8523 7149
rect 5375 6564 8523 6570
rect 5375 6418 8523 6424
rect 5375 5873 5385 6418
rect 5515 6323 6707 6329
rect 7171 6323 8413 6329
rect 5515 6289 5527 6323
rect 6695 6289 7183 6323
rect 8351 6289 8413 6323
rect 5515 6283 6707 6289
rect 7171 6283 8413 6289
rect 8379 6251 8413 6283
rect 5459 6239 5505 6251
rect 5459 6127 5465 6239
rect 5499 6127 5505 6239
rect 6717 6239 6763 6251
rect 6717 6163 6723 6239
rect 6757 6163 6763 6239
rect 7115 6239 7161 6251
rect 8373 6239 8419 6251
rect 7115 6163 7121 6239
rect 7155 6163 7161 6239
rect 8354 6175 8364 6239
rect 8428 6175 8438 6239
rect 5440 6063 5450 6127
rect 5514 6063 5524 6127
rect 6704 6063 6714 6163
rect 6766 6063 6776 6163
rect 7102 6063 7112 6163
rect 7164 6063 7174 6163
rect 8373 6063 8379 6175
rect 8413 6063 8419 6175
rect 5459 6051 5505 6063
rect 6717 6051 6763 6063
rect 7115 6051 7161 6063
rect 8373 6051 8419 6063
rect 8379 6019 8413 6051
rect 5515 6013 6707 6019
rect 7171 6013 8413 6019
rect 5515 5979 5527 6013
rect 6695 5979 7183 6013
rect 8351 5979 8413 6013
rect 5515 5973 6707 5979
rect 7171 5973 8413 5979
rect 8513 5873 8523 6418
rect 5375 5867 8523 5873
rect 5289 5727 5335 5730
rect 5289 5721 8523 5727
rect 5289 5718 5381 5721
rect 8513 5720 8523 5721
rect 8589 5720 8599 7927
rect 8517 5708 8595 5720
rect 13745 2263 13753 11032
rect 20417 10853 20429 11042
rect 13873 10847 16576 10853
rect 13873 2397 13879 10847
rect 14153 10691 14409 10697
rect 14745 10691 15031 10697
rect 15334 10691 15620 10697
rect 15917 10691 16203 10697
rect 14107 10679 14453 10691
rect 14107 10282 14113 10679
rect 14151 10282 14409 10679
rect 14447 10282 14453 10679
rect 14107 10270 14453 10282
rect 14699 10679 15045 10691
rect 14699 10282 14705 10679
rect 14743 10282 15001 10679
rect 15039 10282 15045 10679
rect 14699 10270 15045 10282
rect 15291 10679 15637 10691
rect 15291 10282 15297 10679
rect 15335 10282 15593 10679
rect 15631 10282 15637 10679
rect 15291 10270 15637 10282
rect 15883 10679 16229 10691
rect 15883 10282 15889 10679
rect 15927 10282 16185 10679
rect 16223 10282 16229 10679
rect 15883 10270 16229 10282
rect 14153 10265 14409 10270
rect 14745 10265 15031 10270
rect 15334 10265 15620 10270
rect 15917 10265 16203 10270
rect 16566 9935 16576 10847
rect 20413 10847 20429 10853
rect 16603 9760 20125 9766
rect 16603 9726 16671 9760
rect 16739 9726 16829 9760
rect 16897 9726 16987 9760
rect 17055 9726 17145 9760
rect 17213 9726 17303 9760
rect 17371 9726 17461 9760
rect 17529 9726 17619 9760
rect 17687 9726 17777 9760
rect 17845 9726 17935 9760
rect 18003 9726 18093 9760
rect 18161 9726 18251 9760
rect 18319 9726 18409 9760
rect 18477 9726 18567 9760
rect 18635 9726 18725 9760
rect 18793 9726 18883 9760
rect 18951 9726 19041 9760
rect 19109 9726 19199 9760
rect 19267 9726 19357 9760
rect 19425 9726 19515 9760
rect 19583 9726 19673 9760
rect 19741 9726 19831 9760
rect 19899 9726 19989 9760
rect 20057 9726 20125 9760
rect 16603 9720 20125 9726
rect 16603 9676 16649 9720
rect 16761 9676 16807 9688
rect 16919 9676 16965 9720
rect 17077 9676 17123 9688
rect 17235 9676 17281 9720
rect 17393 9676 17439 9688
rect 17551 9676 17597 9720
rect 17709 9676 17755 9688
rect 17867 9676 17913 9720
rect 18025 9677 18071 9688
rect 16603 8100 16609 9676
rect 16643 8100 16649 9676
rect 16748 9276 16758 9676
rect 16810 9276 16820 9676
rect 16590 7700 16600 8100
rect 16652 7700 16662 8100
rect 16761 7700 16767 9276
rect 16801 7700 16807 9276
rect 16919 8100 16925 9676
rect 16959 8100 16965 9676
rect 17064 9276 17074 9676
rect 17126 9276 17136 9676
rect 16906 7700 16916 8100
rect 16968 7700 16978 8100
rect 17077 7700 17083 9276
rect 17117 7700 17123 9276
rect 17235 8100 17241 9676
rect 17275 8100 17281 9676
rect 17380 9276 17390 9676
rect 17442 9276 17452 9676
rect 17222 7700 17232 8100
rect 17284 7700 17294 8100
rect 17393 7700 17399 9276
rect 17433 7700 17439 9276
rect 17551 8100 17557 9676
rect 17591 8100 17597 9676
rect 17696 9276 17706 9676
rect 17758 9276 17768 9676
rect 17538 7700 17548 8100
rect 17600 7700 17610 8100
rect 17709 7700 17715 9276
rect 17749 7700 17755 9276
rect 17867 8100 17873 9676
rect 17907 8100 17913 9676
rect 18012 9277 18022 9677
rect 18074 9277 18084 9677
rect 18183 9676 18229 9720
rect 18341 9676 18387 9688
rect 18499 9676 18545 9720
rect 18657 9676 18703 9688
rect 18815 9676 18861 9720
rect 18973 9676 19019 9688
rect 19131 9676 19177 9720
rect 19289 9676 19335 9688
rect 19447 9676 19493 9720
rect 19605 9676 19651 9688
rect 19763 9676 19809 9720
rect 19921 9676 19967 9688
rect 20079 9676 20125 9720
rect 17854 7700 17864 8100
rect 17916 7700 17926 8100
rect 18025 7700 18031 9277
rect 18065 7700 18071 9277
rect 18183 8100 18189 9676
rect 18223 8100 18229 9676
rect 18328 9276 18338 9676
rect 18390 9276 18400 9676
rect 18170 7700 18180 8100
rect 18232 7700 18242 8100
rect 18341 7700 18347 9276
rect 18381 7700 18387 9276
rect 18499 8100 18505 9676
rect 18539 8100 18545 9676
rect 18644 9276 18654 9676
rect 18706 9276 18716 9676
rect 18486 7700 18496 8100
rect 18548 7700 18558 8100
rect 18657 7700 18663 9276
rect 18697 7700 18703 9276
rect 18815 8100 18821 9676
rect 18855 8100 18861 9676
rect 18960 9276 18970 9676
rect 19022 9276 19032 9676
rect 18802 7700 18812 8100
rect 18864 7700 18874 8100
rect 18973 7700 18979 9276
rect 19013 7700 19019 9276
rect 19131 8100 19137 9676
rect 19171 8100 19177 9676
rect 19276 9276 19286 9676
rect 19338 9276 19348 9676
rect 19118 7700 19128 8100
rect 19180 7700 19190 8100
rect 19289 7700 19295 9276
rect 19329 7700 19335 9276
rect 19447 8100 19453 9676
rect 19487 8100 19493 9676
rect 19592 9276 19602 9676
rect 19654 9276 19664 9676
rect 19434 7700 19444 8100
rect 19496 7700 19506 8100
rect 19605 7700 19611 9276
rect 19645 7700 19651 9276
rect 19763 8100 19769 9676
rect 19803 8100 19809 9676
rect 19908 9276 19918 9676
rect 19970 9276 19980 9676
rect 19750 7700 19760 8100
rect 19812 7700 19822 8100
rect 19921 7700 19927 9276
rect 19961 7700 19967 9276
rect 20079 8100 20085 9676
rect 20119 8100 20125 9676
rect 20268 9488 20274 9935
rect 20413 9737 20423 10847
rect 20066 7700 20076 8100
rect 20128 7700 20138 8100
rect 16603 7656 16649 7700
rect 16761 7688 16807 7700
rect 16919 7656 16965 7700
rect 17077 7688 17123 7700
rect 17235 7656 17281 7700
rect 17393 7688 17439 7700
rect 17551 7656 17597 7700
rect 17709 7688 17755 7700
rect 17867 7656 17913 7700
rect 18025 7688 18071 7700
rect 18183 7656 18229 7700
rect 18341 7688 18387 7700
rect 18499 7656 18545 7700
rect 18657 7688 18703 7700
rect 18815 7656 18861 7700
rect 18973 7688 19019 7700
rect 19131 7656 19177 7700
rect 19289 7688 19335 7700
rect 19447 7656 19493 7700
rect 19605 7688 19651 7700
rect 19763 7656 19809 7700
rect 19921 7688 19967 7700
rect 20079 7656 20125 7700
rect 16603 7650 20125 7656
rect 16603 7616 16671 7650
rect 16739 7616 16829 7650
rect 16897 7616 16987 7650
rect 17055 7616 17145 7650
rect 17213 7616 17303 7650
rect 17371 7616 17461 7650
rect 17529 7616 17619 7650
rect 17687 7616 17777 7650
rect 17845 7616 17935 7650
rect 18003 7616 18093 7650
rect 18161 7616 18251 7650
rect 18319 7616 18409 7650
rect 18477 7616 18567 7650
rect 18635 7616 18725 7650
rect 18793 7616 18883 7650
rect 18951 7616 19041 7650
rect 19109 7616 19199 7650
rect 19267 7616 19357 7650
rect 19425 7616 19515 7650
rect 19583 7616 19673 7650
rect 19741 7616 19831 7650
rect 19899 7616 19989 7650
rect 20057 7616 20125 7650
rect 16603 7610 20125 7616
rect 20251 7485 20261 9488
rect 20154 7479 20261 7485
rect 16459 7473 20261 7479
rect 16459 7290 16471 7473
rect 16459 7284 18343 7290
rect 18333 7243 18343 7284
rect 14437 7192 14723 7197
rect 15030 7192 15316 7197
rect 15614 7192 15900 7197
rect 14107 7180 14157 7192
rect 14107 6798 14113 7180
rect 14097 6783 14113 6798
rect 14151 6798 14157 7180
rect 14403 7180 14749 7192
rect 14151 6783 14167 6798
rect 14097 6521 14167 6783
rect 14403 6783 14409 7180
rect 14447 6783 14705 7180
rect 14743 6783 14749 7180
rect 14403 6771 14749 6783
rect 14995 7180 15341 7192
rect 14995 6783 15001 7180
rect 15039 6783 15297 7180
rect 15335 6783 15341 7180
rect 14995 6771 15341 6783
rect 15587 7180 15933 7192
rect 16179 7183 16229 7192
rect 16683 7183 16693 7186
rect 15587 6783 15593 7180
rect 15631 6783 15889 7180
rect 15927 6783 15933 7180
rect 16168 6783 16178 7183
rect 16230 6783 16240 7183
rect 16681 7137 16693 7183
rect 16869 7183 16879 7186
rect 17269 7183 17279 7186
rect 16683 7134 16693 7137
rect 16869 7137 16881 7183
rect 17267 7137 17279 7183
rect 17455 7183 17465 7186
rect 17855 7183 17865 7186
rect 16869 7134 16879 7137
rect 17269 7134 17279 7137
rect 17455 7137 17467 7183
rect 17853 7137 17865 7183
rect 18041 7183 18051 7186
rect 17455 7134 17465 7137
rect 17855 7134 17865 7137
rect 18041 7137 18053 7183
rect 18041 7134 18051 7137
rect 16603 7115 16649 7127
rect 15587 6771 15933 6783
rect 16179 6771 16229 6783
rect 14437 6765 14723 6771
rect 15030 6765 15316 6771
rect 15614 6765 15900 6771
rect 14432 6533 14708 6539
rect 15034 6533 15310 6539
rect 15623 6533 15899 6539
rect 14097 6499 14113 6521
rect 14107 6124 14113 6499
rect 14151 6499 14167 6521
rect 14403 6521 14749 6533
rect 14151 6124 14157 6499
rect 14107 6112 14157 6124
rect 14403 6124 14409 6521
rect 14447 6124 14705 6521
rect 14743 6124 14749 6521
rect 14403 6112 14749 6124
rect 14995 6521 15341 6533
rect 14995 6124 15001 6521
rect 15039 6124 15297 6521
rect 15335 6124 15341 6521
rect 14995 6112 15341 6124
rect 15587 6521 15933 6533
rect 15587 6124 15593 6521
rect 15631 6124 15889 6521
rect 15927 6124 15933 6521
rect 15587 6112 15933 6124
rect 14432 6107 14708 6112
rect 15034 6107 15310 6112
rect 15623 6107 15899 6112
rect 16159 6107 16169 6539
rect 16239 6107 16249 6539
rect 16179 6106 16229 6107
rect 16603 5147 16609 7115
rect 16643 7042 16649 7115
rect 16913 7115 17235 7127
rect 16913 7042 16919 7115
rect 16643 5222 16919 7042
rect 16643 5147 16649 5222
rect 16603 5135 16649 5147
rect 16913 5147 16919 5222
rect 16953 5147 17195 7115
rect 17229 7042 17235 7115
rect 17499 7124 17554 7127
rect 17766 7124 17821 7127
rect 17499 7121 17555 7124
rect 17764 7121 17821 7124
rect 17499 7115 17821 7121
rect 17499 7042 17505 7115
rect 17229 5232 17505 7042
rect 17229 5147 17235 5232
rect 16913 5135 17235 5147
rect 17499 5147 17505 5232
rect 17539 5149 17781 7115
rect 17539 5147 17555 5149
rect 17499 5138 17555 5147
rect 17764 5147 17781 5149
rect 17815 7042 17821 7115
rect 18085 7115 18131 7127
rect 18085 7042 18091 7115
rect 17815 5657 18091 7042
rect 18125 5657 18131 7115
rect 18507 6561 19538 6567
rect 18507 6378 18519 6561
rect 19526 6378 19538 6561
rect 18507 6372 19538 6378
rect 18747 6233 19057 6234
rect 19343 6233 19653 6239
rect 18724 6221 19080 6233
rect 18724 5824 18730 6221
rect 18768 5824 19026 6221
rect 19064 5824 19080 6221
rect 18724 5812 19080 5824
rect 19306 6221 19683 6233
rect 19306 5824 19322 6221
rect 19360 5824 19618 6221
rect 19656 5824 19683 6221
rect 19306 5812 19683 5824
rect 18747 5807 19057 5812
rect 17815 5232 18082 5657
rect 17815 5147 17821 5232
rect 18072 5147 18082 5232
rect 18134 5147 18144 5657
rect 17764 5138 17821 5147
rect 17499 5135 17554 5138
rect 17766 5135 17821 5138
rect 18085 5135 18131 5147
rect 16683 5125 16693 5128
rect 16681 5079 16693 5125
rect 16869 5125 16879 5128
rect 17269 5125 17279 5128
rect 16683 5076 16693 5079
rect 16869 5079 16881 5125
rect 17267 5079 17279 5125
rect 17455 5125 17465 5128
rect 17855 5125 17865 5128
rect 16869 5076 16879 5079
rect 17269 5076 17279 5079
rect 17455 5079 17467 5125
rect 17853 5079 17865 5125
rect 18041 5125 18051 5128
rect 17455 5076 17465 5079
rect 17855 5076 17865 5079
rect 18041 5079 18053 5125
rect 18041 5076 18051 5079
rect 16683 4721 16693 4724
rect 16681 4675 16693 4721
rect 16869 4721 16879 4724
rect 17269 4721 17279 4724
rect 16683 4672 16693 4675
rect 16869 4675 16881 4721
rect 17267 4675 17279 4721
rect 17455 4721 17465 4724
rect 17855 4721 17865 4724
rect 16869 4672 16879 4675
rect 17269 4672 17279 4675
rect 17455 4675 17467 4721
rect 17853 4675 17865 4721
rect 18041 4721 18051 4724
rect 17455 4672 17465 4675
rect 17855 4672 17865 4675
rect 18041 4675 18053 4721
rect 18041 4672 18051 4675
rect 16603 4653 16649 4665
rect 14141 3034 14417 3039
rect 14740 3034 15016 3039
rect 15323 3034 15599 3039
rect 15924 3034 16200 3039
rect 14107 3022 14453 3034
rect 14107 2625 14113 3022
rect 14151 2625 14409 3022
rect 14447 2625 14453 3022
rect 14107 2613 14453 2625
rect 14699 3022 15045 3034
rect 14699 2625 14705 3022
rect 14743 2625 15001 3022
rect 15039 2625 15045 3022
rect 14699 2613 15045 2625
rect 15291 3022 15637 3034
rect 15291 2625 15297 3022
rect 15335 2625 15593 3022
rect 15631 2625 15637 3022
rect 15291 2613 15637 2625
rect 15883 3022 16229 3034
rect 15883 2625 15889 3022
rect 15927 2625 16185 3022
rect 16223 2625 16229 3022
rect 16603 2685 16609 4653
rect 16643 2685 16649 4653
rect 16603 2673 16649 2685
rect 16913 4653 17235 4665
rect 16913 2685 16919 4653
rect 16953 2685 17195 4653
rect 17229 2685 17235 4653
rect 16913 2673 17235 2685
rect 17499 4653 17821 4665
rect 17499 2685 17505 4653
rect 17539 2685 17781 4653
rect 17815 2685 17821 4653
rect 18085 4653 18131 4665
rect 18085 3185 18091 4653
rect 18125 3185 18131 4653
rect 18072 2685 18082 3185
rect 18134 2685 18144 3185
rect 17499 2673 17821 2685
rect 18085 2673 18131 2685
rect 16683 2663 16693 2666
rect 15883 2613 16229 2625
rect 16681 2617 16693 2663
rect 16869 2663 16879 2666
rect 17269 2663 17279 2666
rect 16683 2614 16693 2617
rect 16869 2617 16881 2663
rect 17267 2617 17279 2663
rect 17455 2663 17465 2666
rect 17855 2663 17865 2666
rect 16869 2614 16879 2617
rect 17269 2614 17279 2617
rect 17455 2617 17467 2663
rect 17853 2617 17865 2663
rect 18041 2663 18051 2666
rect 17455 2614 17465 2617
rect 17855 2614 17865 2617
rect 18041 2617 18053 2663
rect 18041 2614 18051 2617
rect 14141 2607 14417 2613
rect 14740 2607 15016 2613
rect 15323 2607 15599 2613
rect 15924 2607 16200 2613
rect 18704 2607 18714 3039
rect 18784 2607 18794 3039
rect 19010 3022 19376 3034
rect 19010 2625 19026 3022
rect 19064 2625 19322 3022
rect 19360 2625 19376 3022
rect 19010 2613 19376 2625
rect 19053 2607 19363 2613
rect 19592 2607 19602 3039
rect 19673 2607 19683 3039
rect 20089 2397 20099 7243
rect 13873 2391 20099 2397
rect 13747 2259 13753 2263
rect 13747 2254 20160 2259
rect 20400 2254 20406 9737
rect 24357 8174 24625 8180
rect 24357 8168 25891 8174
rect 21313 8164 24037 8167
rect 21310 8157 21320 8164
rect 21189 8145 21320 8157
rect 21185 3233 21195 8145
rect 24092 8022 24102 8164
rect 21504 5970 21514 8022
rect 22995 7951 23005 7954
rect 21737 7945 23005 7951
rect 23725 7951 23735 7954
rect 21737 7911 21749 7945
rect 21737 7905 23005 7911
rect 22995 7902 23005 7905
rect 23725 7905 23737 7951
rect 23725 7902 23735 7905
rect 21659 7883 21705 7895
rect 21659 7127 21665 7883
rect 21699 7809 21705 7883
rect 23769 7883 23815 7895
rect 23769 7809 23775 7883
rect 21699 7127 23775 7809
rect 21644 6127 21654 7127
rect 21710 6189 23775 7127
rect 21710 6127 21720 6189
rect 21659 6115 21665 6127
rect 21699 6115 21705 6127
rect 21659 6103 21705 6115
rect 23767 6115 23775 6189
rect 23809 6712 23815 7883
rect 23905 7809 23911 8022
rect 24090 7809 24096 8022
rect 24357 7835 24363 8168
rect 25879 8165 25891 8168
rect 25879 8161 26801 8165
rect 25879 8159 26841 8161
rect 24619 8034 25836 8040
rect 24619 7835 24625 8034
rect 24357 7823 24364 7835
rect 23809 6115 23834 6712
rect 21739 6093 21749 6096
rect 21737 6047 21749 6093
rect 22469 6093 22479 6096
rect 22469 6087 23737 6093
rect 23725 6053 23737 6087
rect 21739 6044 21749 6047
rect 22469 6047 23737 6053
rect 22469 6044 22479 6047
rect 21504 5964 23735 5970
rect 23723 5795 23735 5964
rect 23767 5837 23834 6115
rect 21504 5789 23735 5795
rect 21504 3597 21514 5789
rect 21659 5787 21705 5789
rect 21739 5701 21749 5704
rect 21737 5655 21749 5701
rect 22469 5701 22479 5704
rect 22469 5695 23737 5701
rect 23725 5661 23737 5695
rect 21739 5652 21749 5655
rect 22469 5655 23737 5661
rect 22469 5652 22479 5655
rect 21659 5633 21705 5650
rect 21659 5608 21665 5633
rect 21699 5608 21705 5633
rect 23766 5633 23834 5837
rect 21644 5285 21654 5608
rect 21710 5544 21720 5608
rect 23766 5544 23775 5633
rect 21710 5285 23775 5544
rect 21659 4865 21665 5285
rect 21699 4865 23775 5285
rect 21643 3865 21653 4865
rect 21709 3943 23775 4865
rect 21709 3865 21719 3943
rect 23769 3865 23775 3943
rect 23809 5436 23834 5633
rect 23809 5191 23833 5436
rect 23809 3930 23815 5191
rect 23899 4053 23909 7809
rect 24092 4317 24102 7809
rect 24358 7772 24364 7823
rect 24618 7823 24625 7835
rect 24744 7902 24843 7954
rect 25413 7951 25423 7954
rect 25413 7945 25718 7951
rect 25619 7911 25718 7945
rect 25413 7905 25718 7911
rect 25413 7902 25423 7905
rect 24744 7883 24790 7902
rect 24618 7772 24624 7823
rect 24354 5031 24364 7772
rect 24346 5025 24364 5031
rect 24618 5031 24628 7772
rect 24744 7715 24750 7883
rect 24784 7855 24790 7883
rect 25672 7883 25718 7905
rect 25672 7855 25678 7883
rect 24784 7730 25678 7855
rect 24784 7715 24790 7730
rect 24744 7177 24790 7715
rect 25672 7715 25678 7730
rect 25712 7715 25718 7883
rect 25672 7703 25718 7715
rect 25039 7693 25049 7696
rect 24831 7687 25049 7693
rect 25619 7693 25629 7696
rect 24831 7653 24843 7687
rect 24831 7647 25049 7653
rect 25039 7644 25049 7647
rect 25619 7647 25631 7693
rect 25619 7644 25629 7647
rect 25824 7543 25836 8034
rect 24871 7537 25836 7543
rect 24871 7354 24883 7537
rect 25918 7363 26708 7369
rect 25918 7354 25930 7363
rect 24871 7348 25930 7354
rect 24833 7245 24843 7248
rect 24831 7199 24843 7245
rect 25563 7245 25573 7248
rect 25563 7239 26531 7245
rect 26519 7205 26531 7239
rect 24833 7196 24843 7199
rect 25563 7199 26531 7205
rect 25563 7196 25573 7199
rect 24744 7009 24750 7177
rect 24784 7009 24790 7177
rect 24744 6919 24790 7009
rect 26572 7177 26618 7193
rect 26572 7009 26578 7177
rect 26612 7009 26618 7177
rect 25789 6987 25799 6990
rect 24831 6981 25799 6987
rect 26519 6987 26529 6990
rect 24831 6947 24843 6981
rect 24831 6941 25799 6947
rect 25789 6938 25799 6941
rect 26519 6941 26531 6987
rect 26519 6938 26529 6941
rect 24744 6751 24750 6919
rect 24784 6751 24790 6919
rect 24744 6661 24790 6751
rect 26572 6919 26618 7009
rect 26572 6751 26578 6919
rect 26612 6751 26618 6919
rect 24833 6729 24843 6732
rect 24831 6683 24843 6729
rect 25563 6729 25573 6732
rect 25563 6723 26531 6729
rect 26519 6689 26531 6723
rect 24833 6680 24843 6683
rect 25563 6683 26531 6689
rect 25563 6680 25573 6683
rect 24744 6493 24750 6661
rect 24784 6493 24790 6661
rect 24744 6403 24790 6493
rect 26572 6661 26618 6751
rect 26572 6493 26578 6661
rect 26612 6493 26618 6661
rect 25789 6471 25799 6474
rect 24831 6465 25799 6471
rect 26519 6471 26529 6474
rect 24831 6431 24843 6465
rect 24831 6425 25799 6431
rect 25789 6422 25799 6425
rect 26519 6425 26531 6471
rect 26519 6422 26529 6425
rect 24744 6235 24750 6403
rect 24784 6235 24790 6403
rect 24744 6145 24790 6235
rect 26572 6403 26618 6493
rect 26572 6235 26578 6403
rect 26612 6235 26618 6403
rect 24833 6213 24843 6216
rect 24831 6167 24843 6213
rect 25563 6213 25573 6216
rect 25563 6207 26531 6213
rect 26519 6173 26531 6207
rect 24833 6164 24843 6167
rect 25563 6167 26531 6173
rect 25563 6164 25573 6167
rect 24744 5977 24750 6145
rect 24784 5977 24790 6145
rect 24744 5887 24790 5977
rect 26572 6145 26618 6235
rect 26572 5977 26578 6145
rect 26612 5977 26618 6145
rect 25789 5955 25799 5958
rect 24831 5949 25799 5955
rect 26519 5955 26529 5958
rect 24831 5915 24843 5949
rect 24831 5909 25799 5915
rect 25789 5906 25799 5909
rect 26519 5909 26531 5955
rect 26519 5906 26529 5909
rect 24744 5719 24750 5887
rect 24784 5719 24790 5887
rect 24744 5629 24790 5719
rect 26572 5887 26618 5977
rect 26572 5719 26578 5887
rect 26612 5719 26618 5887
rect 24833 5697 24843 5700
rect 24831 5651 24843 5697
rect 25563 5697 25573 5700
rect 25563 5691 26531 5697
rect 26519 5657 26531 5691
rect 24833 5648 24843 5651
rect 25563 5651 26531 5657
rect 25563 5648 25573 5651
rect 24744 5461 24750 5629
rect 24784 5461 24790 5629
rect 24744 5371 24790 5461
rect 26572 5629 26618 5719
rect 26572 5461 26578 5629
rect 26612 5461 26618 5629
rect 26698 5601 26708 7363
rect 26835 5601 26845 8159
rect 25790 5439 25800 5442
rect 24831 5433 25800 5439
rect 26520 5439 26530 5442
rect 24831 5399 24843 5433
rect 24831 5393 25800 5399
rect 25790 5390 25800 5393
rect 26520 5393 26531 5439
rect 26520 5390 26530 5393
rect 26572 5371 26618 5461
rect 24729 5203 24739 5371
rect 24795 5203 24805 5371
rect 26572 5203 26578 5371
rect 26612 5203 26618 5371
rect 26702 5334 26708 5601
rect 26835 5334 26841 5601
rect 24744 5191 24790 5203
rect 26572 5191 26618 5203
rect 24833 5181 24843 5184
rect 24831 5135 24843 5181
rect 25563 5181 25573 5184
rect 25563 5175 26531 5181
rect 26519 5141 26531 5175
rect 24833 5132 24843 5135
rect 25563 5135 26531 5141
rect 25563 5132 25573 5135
rect 26699 5031 26708 5334
rect 24618 5025 26708 5031
rect 24346 4469 24358 5025
rect 26836 4535 26846 5334
rect 26836 4492 26847 4535
rect 26835 4469 26847 4492
rect 24346 4463 26847 4469
rect 26824 4317 26911 4323
rect 24092 4311 26917 4317
rect 23905 4050 24020 4053
rect 23905 4047 26830 4050
rect 24008 4044 26830 4047
rect 23809 3865 23816 3930
rect 21659 3853 21705 3865
rect 23769 3859 23816 3865
rect 23769 3853 23815 3859
rect 22995 3843 23005 3846
rect 21737 3837 23005 3843
rect 23725 3843 23735 3846
rect 24668 3843 24678 3846
rect 21737 3803 21749 3837
rect 21737 3797 23005 3803
rect 22995 3794 23005 3797
rect 23725 3797 23737 3843
rect 24666 3797 24678 3843
rect 25398 3843 25408 3846
rect 25398 3837 26666 3843
rect 26654 3803 26666 3837
rect 23725 3794 23735 3797
rect 24668 3794 24678 3797
rect 25398 3797 26666 3803
rect 25398 3794 25408 3797
rect 24588 3775 24634 3787
rect 23905 3744 24096 3756
rect 23905 3597 23911 3744
rect 21504 3591 23911 3597
rect 24090 3597 24096 3744
rect 24588 3715 24594 3775
rect 24628 3715 24634 3775
rect 26698 3775 26744 3787
rect 24090 3591 24313 3597
rect 24301 3274 24313 3591
rect 24301 3246 24325 3274
rect 21187 3100 21199 3233
rect 24301 3201 24313 3246
rect 24295 3195 24313 3201
rect 21193 2403 21199 3100
rect 21328 3100 24187 3106
rect 21328 2403 21334 3100
rect 21496 2999 24010 3005
rect 21496 2965 21508 2999
rect 21676 2965 21766 2999
rect 21934 2965 22024 2999
rect 22192 2965 22282 2999
rect 22450 2965 22540 2999
rect 22708 2965 22798 2999
rect 22966 2965 23056 2999
rect 23224 2965 23314 2999
rect 23482 2965 23572 2999
rect 23740 2965 23830 2999
rect 23998 2965 24010 2999
rect 21496 2959 24010 2965
rect 21440 2915 21486 2927
rect 21427 2715 21437 2915
rect 21489 2715 21499 2915
rect 13747 2253 20406 2254
rect 13747 2247 13879 2253
rect 18624 2249 18674 2253
rect 20154 2242 20406 2253
rect 21013 2035 21023 2403
rect 21328 2035 21338 2403
rect 21193 1656 21199 2035
rect 21328 1790 21334 2035
rect 21440 1939 21446 2715
rect 21480 1939 21486 2715
rect 21440 1927 21486 1939
rect 21533 1898 21650 2959
rect 21698 2915 21744 2927
rect 21698 2139 21704 2915
rect 21738 2139 21744 2915
rect 21685 1939 21695 2139
rect 21747 1939 21757 2139
rect 21698 1927 21744 1939
rect 21498 1895 21508 1898
rect 21496 1849 21508 1895
rect 21639 1895 21650 1898
rect 21798 1895 21915 2959
rect 21956 2915 22002 2927
rect 21943 2715 21953 2915
rect 22005 2715 22015 2915
rect 21956 1939 21962 2715
rect 21996 1939 22002 2715
rect 21956 1927 22002 1939
rect 22054 1895 22171 2959
rect 22214 2915 22260 2927
rect 22214 2139 22220 2915
rect 22254 2139 22260 2915
rect 22201 1939 22211 2139
rect 22263 1939 22273 2139
rect 22214 1927 22260 1939
rect 22314 1895 22431 2959
rect 22472 2915 22518 2927
rect 22459 2715 22469 2915
rect 22521 2715 22531 2915
rect 22472 1939 22478 2715
rect 22512 1939 22518 2715
rect 22472 1927 22518 1939
rect 22562 1895 22679 2959
rect 22730 2915 22776 2927
rect 22730 2139 22736 2915
rect 22770 2139 22776 2915
rect 22717 1939 22727 2139
rect 22779 1939 22789 2139
rect 22730 1927 22776 1939
rect 22827 1895 22944 2959
rect 22988 2915 23034 2927
rect 22975 2715 22985 2915
rect 23037 2715 23047 2915
rect 22988 1939 22994 2715
rect 23028 1939 23034 2715
rect 22988 1927 23034 1939
rect 23081 1895 23198 2959
rect 23246 2915 23292 2927
rect 23246 2139 23252 2915
rect 23286 2139 23292 2915
rect 23233 1939 23243 2139
rect 23295 1939 23305 2139
rect 23246 1927 23292 1939
rect 23343 1895 23460 2959
rect 23504 2915 23550 2927
rect 23491 2715 23501 2915
rect 23553 2715 23563 2915
rect 23504 1939 23510 2715
rect 23544 1939 23550 2715
rect 23504 1927 23550 1939
rect 23603 1895 23720 2959
rect 23762 2915 23808 2927
rect 23762 2139 23768 2915
rect 23802 2139 23808 2915
rect 23749 1939 23759 2139
rect 23811 1939 23821 2139
rect 23762 1927 23808 1939
rect 23860 1895 23977 2959
rect 24020 2915 24066 2927
rect 24007 2715 24017 2915
rect 24069 2715 24079 2915
rect 24020 1939 24026 2715
rect 24060 1939 24066 2715
rect 24020 1927 24066 1939
rect 21639 1889 24010 1895
rect 21676 1855 21766 1889
rect 21934 1855 22024 1889
rect 22192 1855 22282 1889
rect 22450 1855 22540 1889
rect 22708 1855 22798 1889
rect 22966 1855 23056 1889
rect 23224 1855 23314 1889
rect 23482 1855 23572 1889
rect 23740 1855 23830 1889
rect 23998 1855 24010 1889
rect 21498 1846 21508 1849
rect 21639 1849 24010 1855
rect 21639 1846 21650 1849
rect 24177 1790 24187 3100
rect 21328 1784 24187 1790
rect 24295 1860 24305 3195
rect 24568 2815 24578 3715
rect 24642 3668 24652 3715
rect 26698 3668 26704 3775
rect 24642 2815 26704 3668
rect 24588 2007 24594 2815
rect 24628 2089 26704 2815
rect 24628 2007 24634 2089
rect 26632 2088 26704 2089
rect 24588 1995 24634 2007
rect 26698 2007 26704 2088
rect 26738 2007 26744 3775
rect 26698 1995 26744 2007
rect 24668 1985 24678 1987
rect 24666 1939 24678 1985
rect 25398 1985 25408 1987
rect 25398 1979 26666 1985
rect 26654 1945 26666 1979
rect 24668 1935 24678 1939
rect 25398 1939 26666 1945
rect 25398 1935 25408 1939
rect 26820 1860 26830 4044
rect 24295 1855 26830 1860
rect 24295 1854 26479 1855
rect 26905 4044 26917 4311
rect 26905 1663 26915 4044
rect 24295 1657 26911 1663
rect 24295 1656 24307 1657
rect 21193 1650 24307 1656
rect 21193 1644 21334 1650
<< via1 >>
rect 2433 42577 2669 42578
rect 2669 42577 5829 42578
rect 2433 42347 5829 42577
rect 2433 30250 2681 42347
rect 2681 30250 2688 42347
rect 5603 31000 5613 42347
rect 5613 31000 5815 42347
rect 6032 31118 10883 31303
rect 2784 30763 2856 30766
rect 2784 30366 2802 30763
rect 2802 30366 2840 30763
rect 2840 30366 2856 30763
rect 5459 30366 5466 30763
rect 5466 30366 5504 30763
rect 5504 30366 5511 30763
rect 6224 30730 6233 30830
rect 6233 30730 6267 30830
rect 6267 30730 6276 30830
rect 10602 30806 10617 30906
rect 10617 30806 10651 30906
rect 10651 30806 10666 30906
rect 6295 30671 6548 30679
rect 10229 30671 10589 30686
rect 6295 30637 6548 30671
rect 10229 30637 10589 30671
rect 6295 30622 6548 30637
rect 10229 30613 10589 30637
rect 10759 30536 10874 31118
rect 6031 30351 10882 30536
rect 2429 30063 2431 30250
rect 2431 30245 2681 30250
rect 2681 30245 5613 30250
rect 5613 30245 5815 30250
rect 2431 30063 5815 30245
rect 6236 27582 7095 27983
rect 5742 24614 5981 24621
rect 12861 27801 13258 27808
rect 12861 27763 13258 27801
rect 12861 27756 13258 27763
rect 12958 25137 13258 25144
rect 12958 25099 13258 25137
rect 12958 25092 13258 25099
rect 13986 27792 14066 27818
rect 13986 27758 14031 27792
rect 14031 27758 14065 27792
rect 14065 27758 14066 27792
rect 13986 27692 14066 27758
rect 13986 27658 14031 27692
rect 14031 27658 14065 27692
rect 14065 27658 14066 27692
rect 13986 27592 14066 27658
rect 13986 27558 14031 27592
rect 14031 27558 14065 27592
rect 14065 27558 14066 27592
rect 13986 27492 14066 27558
rect 13986 27458 14031 27492
rect 14031 27458 14065 27492
rect 14065 27458 14066 27492
rect 13986 27392 14066 27458
rect 13986 27358 14031 27392
rect 14031 27358 14065 27392
rect 14065 27358 14066 27392
rect 13986 27344 14066 27358
rect 5742 24599 11232 24614
rect 5742 24211 12844 24599
rect 15378 26048 15907 26070
rect 15378 26014 15409 26048
rect 15409 26014 15475 26048
rect 15475 26014 15509 26048
rect 15509 26014 15575 26048
rect 15575 26014 15609 26048
rect 15609 26014 15675 26048
rect 15675 26014 15709 26048
rect 15709 26014 15775 26048
rect 15775 26014 15809 26048
rect 15809 26014 15875 26048
rect 15875 26014 15907 26048
rect 15378 25984 15907 26014
rect 5742 24198 11232 24211
rect 11232 24204 12844 24211
rect 5742 19777 5981 24198
rect 6180 24068 6240 24102
rect 6180 24050 6240 24068
rect 6280 22961 6290 23961
rect 6290 22961 6324 23961
rect 6324 22961 6332 23961
rect 6180 20044 6240 20050
rect 6180 20010 6240 20044
rect 6180 19998 6240 20010
rect 6650 24068 6710 24102
rect 6650 24050 6710 24068
rect 6558 22961 6566 23961
rect 6566 22961 6600 23961
rect 6600 22961 6610 23961
rect 6768 22961 6776 23961
rect 6776 22961 6810 23961
rect 6810 22961 6820 23961
rect 6666 20010 6726 20044
rect 6666 19992 6726 20010
rect 7152 24102 7212 24120
rect 7152 24068 7212 24102
rect 7046 22963 7052 23963
rect 7052 22963 7086 23963
rect 7086 22963 7098 23963
rect 7136 20010 7196 20044
rect 7136 19992 7196 20010
rect 7638 24102 7698 24120
rect 7638 24068 7698 24102
rect 7737 22966 7748 23966
rect 7748 22966 7782 23966
rect 7782 22966 7789 23966
rect 7622 20010 7682 20044
rect 7622 19992 7682 20010
rect 8108 24102 8168 24120
rect 8108 24068 8168 24102
rect 8016 22966 8024 23966
rect 8024 22966 8058 23966
rect 8058 22966 8068 23966
rect 8225 22964 8234 23964
rect 8234 22964 8268 23964
rect 8268 22964 8277 23964
rect 8124 20010 8184 20044
rect 8124 19992 8184 20010
rect 8610 24102 8670 24120
rect 8610 24068 8670 24102
rect 8500 22964 8510 23964
rect 8510 22964 8544 23964
rect 8544 22964 8552 23964
rect 8712 22963 8720 23963
rect 8720 22963 8754 23963
rect 8754 22963 8764 23963
rect 8594 20010 8654 20044
rect 8594 19992 8654 20010
rect 9080 24102 9140 24120
rect 9080 24068 9140 24102
rect 8987 22963 8996 23963
rect 8996 22963 9030 23963
rect 9030 22963 9039 23963
rect 9197 22963 9206 23963
rect 9206 22963 9240 23963
rect 9240 22963 9249 23963
rect 9096 20010 9156 20044
rect 9096 19992 9156 20010
rect 9582 24102 9642 24120
rect 9582 24068 9642 24102
rect 9473 22963 9482 23963
rect 9482 22963 9516 23963
rect 9516 22963 9525 23963
rect 9684 22963 9692 23963
rect 9692 22963 9726 23963
rect 9726 22963 9736 23963
rect 9566 20010 9626 20044
rect 9566 19992 9626 20010
rect 10052 24102 10112 24120
rect 10052 24068 10112 24102
rect 9959 22963 9968 23963
rect 9968 22963 10002 23963
rect 10002 22963 10011 23963
rect 10169 22963 10178 23963
rect 10178 22963 10212 23963
rect 10212 22963 10221 23963
rect 10068 20010 10128 20044
rect 10068 19992 10128 20010
rect 10554 24102 10614 24120
rect 10554 24068 10614 24102
rect 10446 22963 10454 23963
rect 10454 22963 10488 23963
rect 10488 22963 10498 23963
rect 10538 20010 10598 20044
rect 10538 19992 10598 20010
rect 15564 23789 20117 24049
rect 15788 23407 15797 23607
rect 15797 23407 15831 23607
rect 15831 23407 15840 23607
rect 11332 22631 11341 22831
rect 11341 22631 11375 22831
rect 11375 22631 11384 22831
rect 15390 22631 15399 22831
rect 15399 22631 15433 22831
rect 15433 22631 15442 22831
rect 19846 23407 19855 23607
rect 19855 23407 19889 23607
rect 19889 23407 19898 23607
rect 11352 22172 15126 22356
rect 16147 22146 20041 22381
rect 11339 20959 11348 21159
rect 11348 20959 11382 21159
rect 11382 20959 11391 21159
rect 15530 21187 15686 21768
rect 15788 21735 15797 21935
rect 15797 21735 15831 21935
rect 15831 21735 15840 21935
rect 19846 21735 19855 21935
rect 19855 21735 19889 21935
rect 19889 21735 19898 21935
rect 19961 21189 19965 21752
rect 19965 21189 20148 21752
rect 19961 21187 20148 21189
rect 15530 21161 20148 21187
rect 15397 20959 15406 21159
rect 15406 20959 15440 21159
rect 15440 20959 15449 21159
rect 15537 21110 20148 21161
rect 11279 20696 15029 20783
rect 9350 19132 10350 19143
rect 9350 19098 10350 19132
rect 9350 19087 10350 19098
rect 6349 18763 6358 19039
rect 6358 18763 6392 19039
rect 6392 18763 6401 19039
rect 10407 18763 10416 19039
rect 10416 18763 10450 19039
rect 10450 18763 10459 19039
rect 6349 18227 6358 18503
rect 6358 18227 6392 18503
rect 6392 18227 6401 18503
rect 10407 18227 10416 18503
rect 10416 18227 10450 18503
rect 10450 18227 10459 18503
rect 6342 17439 6358 17639
rect 6358 17439 6392 17639
rect 6392 17439 6406 17639
rect 10407 17063 10416 17639
rect 10416 17063 10450 17639
rect 10450 17063 10459 17639
rect 8420 14928 9420 14937
rect 8420 14894 8430 14928
rect 8430 14894 9420 14928
rect 8420 14885 9420 14894
rect 8054 14450 8056 14789
rect 8056 14464 8243 14789
rect 8243 14464 8246 14789
rect 8349 14659 8368 14786
rect 8368 14659 8401 14786
rect 10407 14659 10416 14835
rect 10416 14659 10450 14835
rect 10450 14659 10459 14835
rect 11506 19132 12506 19143
rect 11506 19098 11508 19132
rect 11508 19098 12506 19132
rect 11506 19087 12506 19098
rect 11431 17063 11446 17663
rect 11446 17063 11480 17663
rect 11480 17063 11495 17663
rect 15495 17063 15504 17563
rect 15504 17063 15538 17563
rect 15538 17063 15547 17563
rect 15763 17063 15772 17563
rect 15772 17063 15806 17563
rect 15806 17063 15815 17563
rect 19815 18439 19830 19039
rect 19830 18439 19864 19039
rect 19864 18439 19879 19039
rect 11431 16035 11446 16635
rect 11446 16035 11480 16635
rect 11480 16035 11495 16635
rect 15495 16135 15504 16635
rect 15504 16135 15538 16635
rect 15538 16135 15547 16635
rect 15763 16135 15772 16635
rect 15772 16135 15806 16635
rect 15806 16135 15815 16635
rect 15495 14659 15504 14850
rect 15504 14659 15538 14850
rect 15538 14659 15547 14850
rect 15763 14659 15772 14850
rect 15772 14659 15806 14850
rect 15806 14659 15815 14850
rect 19815 14792 19830 15259
rect 19830 14792 19864 15259
rect 19864 14792 19879 15259
rect 20911 18768 20987 18780
rect 20911 18734 20987 18768
rect 20911 18728 20987 18734
rect 21403 18768 21503 18796
rect 21403 18734 21415 18768
rect 21415 18734 21491 18768
rect 21491 18734 21503 18768
rect 21403 18732 21503 18734
rect 21035 17700 21046 18700
rect 21046 17700 21080 18700
rect 21080 17700 21091 18700
rect 21539 17658 21550 18658
rect 21550 17658 21584 18658
rect 21584 17658 21595 18658
rect 20911 14710 20987 14716
rect 20911 14676 20987 14710
rect 20911 14664 20987 14676
rect 21415 14710 21491 14716
rect 21415 14676 21491 14710
rect 21415 14664 21491 14676
rect 8056 14454 21806 14464
rect 8056 14418 21822 14454
rect 8056 14001 21806 14418
rect 21806 14001 21822 14418
rect 21564 13991 21822 14001
rect 7800 12663 10778 12824
rect 7800 12519 10779 12663
rect 8064 12311 8116 12335
rect 8064 12135 8073 12311
rect 8073 12135 8107 12311
rect 8107 12135 8116 12311
rect 10122 12135 10141 12311
rect 10141 12135 10174 12311
rect 8135 12076 8844 12084
rect 8135 12042 8844 12076
rect 8135 12032 8844 12042
rect 5836 11194 5840 11969
rect 5840 11761 10075 11969
rect 5840 11194 5983 11761
rect 6058 11172 6073 11548
rect 6073 11172 6107 11548
rect 6107 11172 6116 11548
rect 10122 11172 10131 11548
rect 10131 11172 10165 11548
rect 10165 11172 10174 11548
rect 6135 11113 7135 11115
rect 6135 11079 7135 11113
rect 6135 11063 7135 11079
rect 5840 10840 9712 10956
rect 6170 10327 6185 10562
rect 6185 10327 6219 10562
rect 6219 10327 6234 10562
rect 6892 9970 6985 10194
rect 7644 10086 7659 10322
rect 7659 10086 7693 10322
rect 7693 10086 7708 10322
rect 6235 9818 6335 9918
rect 6607 9668 6707 9768
rect 6170 9044 6185 9280
rect 6185 9044 6219 9280
rect 6219 9044 6234 9280
rect 7171 9818 7271 9918
rect 7549 9668 7649 9768
rect 7644 9285 7659 9520
rect 7659 9285 7693 9520
rect 7693 9285 7708 9520
rect 7787 8871 7942 10840
rect 5870 8767 7960 8871
rect 8812 8863 8950 10840
rect 10284 10806 10779 12519
rect 11880 11114 12899 11117
rect 9036 10104 9051 10304
rect 9051 10104 9085 10304
rect 9085 10104 9100 10304
rect 9580 10380 9589 10580
rect 9589 10380 9623 10580
rect 9623 10380 9632 10580
rect 9974 10380 9983 10580
rect 9983 10380 10017 10580
rect 10017 10380 10026 10580
rect 10506 10380 10521 10580
rect 10521 10380 10555 10580
rect 10555 10380 10570 10580
rect 9036 9295 9051 9495
rect 9051 9295 9085 9495
rect 9085 9295 9100 9495
rect 9580 9295 9589 9495
rect 9589 9295 9623 9495
rect 9623 9295 9632 9495
rect 9974 9295 9983 9495
rect 9983 9295 10017 9495
rect 10017 9295 10026 9495
rect 10506 9019 10521 9219
rect 10521 9019 10555 9219
rect 10555 9019 10570 9219
rect 10655 8863 10776 10806
rect 8812 8741 10776 8863
rect 8821 8737 10776 8741
rect 10655 8728 10776 8737
rect 11848 11079 12899 11114
rect 11848 11006 12901 11079
rect 11848 10404 11967 11006
rect 12024 10677 12033 10777
rect 12033 10677 12067 10777
rect 12067 10677 12076 10777
rect 12340 10753 12349 10853
rect 12349 10753 12383 10853
rect 12383 10753 12392 10853
rect 12656 10677 12665 10777
rect 12665 10677 12699 10777
rect 12699 10677 12708 10777
rect 12148 10295 12203 10349
rect 11241 9287 11310 9898
rect 12330 10172 12384 10226
rect 12773 10418 12901 11006
rect 20291 11032 20413 11040
rect 11408 9558 11417 9638
rect 11417 9558 11451 9638
rect 11451 9558 11460 9638
rect 11566 9462 11575 9542
rect 11575 9462 11609 9542
rect 11609 9462 11618 9542
rect 12122 9558 12131 9638
rect 12131 9558 12165 9638
rect 12165 9558 12174 9638
rect 11964 9462 11973 9542
rect 11973 9462 12007 9542
rect 12007 9462 12016 9542
rect 12035 9378 12103 9412
rect 12035 9356 12103 9378
rect 12520 9558 12529 9638
rect 12529 9558 12563 9638
rect 12563 9558 12572 9638
rect 12678 9462 12687 9542
rect 12687 9462 12721 9542
rect 12721 9462 12730 9542
rect 13234 9558 13243 9638
rect 13243 9558 13277 9638
rect 13277 9558 13286 9638
rect 13076 9462 13085 9542
rect 13085 9462 13119 9542
rect 13119 9462 13128 9542
rect 13147 9378 13215 9412
rect 13147 9356 13215 9378
rect 13384 9287 13448 9900
rect 11241 9173 13446 9287
rect 8523 8640 8589 8650
rect 5318 8630 8589 8640
rect 5295 8626 8589 8630
rect 5295 8564 10790 8626
rect 5295 8560 8589 8564
rect 5295 8009 5375 8560
rect 5450 8323 5465 8387
rect 5465 8323 5499 8387
rect 5499 8323 5514 8387
rect 6714 8287 6723 8387
rect 6723 8287 6757 8387
rect 6757 8287 6766 8387
rect 7112 8287 7121 8387
rect 7121 8287 7155 8387
rect 7155 8287 7164 8387
rect 8364 8211 8379 8275
rect 8379 8211 8413 8275
rect 8413 8211 8428 8275
rect 8523 8009 8589 8560
rect 5295 7995 8589 8009
rect 8824 7995 8961 8564
rect 9036 8287 9051 8387
rect 9051 8287 9085 8387
rect 9085 8287 9100 8387
rect 9540 8211 9549 8311
rect 9549 8211 9583 8311
rect 9583 8211 9592 8311
rect 9113 8161 9273 8171
rect 9113 8127 9273 8161
rect 9113 8107 9273 8127
rect 9704 7995 9897 8564
rect 10014 8288 10023 8388
rect 10023 8288 10057 8388
rect 10057 8288 10066 8388
rect 10506 8288 10521 8388
rect 10521 8288 10555 8388
rect 10555 8288 10570 8388
rect 10085 8162 10245 8173
rect 10085 8128 10245 8162
rect 10085 8109 10245 8128
rect 10665 7995 10790 8564
rect 5295 7933 10802 7995
rect 5295 7869 8589 7933
rect 5295 7295 5375 7869
rect 5450 7607 5465 7671
rect 5465 7607 5499 7671
rect 5499 7607 5514 7671
rect 6714 7495 6723 7595
rect 6723 7495 6757 7595
rect 6757 7495 6766 7595
rect 7112 7495 7121 7595
rect 7121 7495 7155 7595
rect 7155 7495 7164 7595
rect 8364 7495 8379 7548
rect 8379 7495 8413 7548
rect 8413 7495 8428 7548
rect 8364 7484 8428 7495
rect 8523 7295 8589 7869
rect 5295 7155 8589 7295
rect 5295 6564 5375 7155
rect 5450 6891 5465 6955
rect 5465 6891 5499 6955
rect 5499 6891 5514 6955
rect 8364 6891 8379 6955
rect 8379 6891 8413 6955
rect 8413 6891 8428 6955
rect 6714 6779 6723 6879
rect 6723 6779 6757 6879
rect 6757 6779 6766 6879
rect 7112 6779 7121 6879
rect 7121 6779 7155 6879
rect 7155 6779 7164 6879
rect 8523 6564 8589 7155
rect 5295 6424 8589 6564
rect 5295 5867 5375 6424
rect 8364 6175 8379 6239
rect 8379 6175 8413 6239
rect 8413 6175 8428 6239
rect 5450 6063 5465 6127
rect 5465 6063 5499 6127
rect 5499 6063 5514 6127
rect 6714 6063 6723 6163
rect 6723 6063 6757 6163
rect 6757 6063 6766 6163
rect 7112 6063 7121 6163
rect 7121 6063 7155 6163
rect 7155 6063 7164 6163
rect 8523 5867 8589 6424
rect 5295 5730 8589 5867
rect 5335 5727 8589 5730
rect 8523 5720 8589 5727
rect 13755 10864 20413 11032
rect 13755 2384 13869 10864
rect 16576 10853 20413 10864
rect 16576 10288 20413 10853
rect 16576 10100 16585 10288
rect 16585 10277 20388 10288
rect 20388 10277 20413 10288
rect 16585 10100 20400 10277
rect 16576 9935 20274 10100
rect 20274 9935 20400 10100
rect 16758 9276 16767 9676
rect 16767 9276 16801 9676
rect 16801 9276 16810 9676
rect 16600 7700 16609 8100
rect 16609 7700 16643 8100
rect 16643 7700 16652 8100
rect 17074 9276 17083 9676
rect 17083 9276 17117 9676
rect 17117 9276 17126 9676
rect 16916 7700 16925 8100
rect 16925 7700 16959 8100
rect 16959 7700 16968 8100
rect 17390 9276 17399 9676
rect 17399 9276 17433 9676
rect 17433 9276 17442 9676
rect 17232 7700 17241 8100
rect 17241 7700 17275 8100
rect 17275 7700 17284 8100
rect 17706 9276 17715 9676
rect 17715 9276 17749 9676
rect 17749 9276 17758 9676
rect 17548 7700 17557 8100
rect 17557 7700 17591 8100
rect 17591 7700 17600 8100
rect 18022 9676 18074 9677
rect 18022 9277 18031 9676
rect 18031 9277 18065 9676
rect 18065 9277 18074 9676
rect 17864 7700 17873 8100
rect 17873 7700 17907 8100
rect 17907 7700 17916 8100
rect 18338 9276 18347 9676
rect 18347 9276 18381 9676
rect 18381 9276 18390 9676
rect 18180 7700 18189 8100
rect 18189 7700 18223 8100
rect 18223 7700 18232 8100
rect 18654 9276 18663 9676
rect 18663 9276 18697 9676
rect 18697 9276 18706 9676
rect 18496 7700 18505 8100
rect 18505 7700 18539 8100
rect 18539 7700 18548 8100
rect 18970 9276 18979 9676
rect 18979 9276 19013 9676
rect 19013 9276 19022 9676
rect 18812 7700 18821 8100
rect 18821 7700 18855 8100
rect 18855 7700 18864 8100
rect 19286 9276 19295 9676
rect 19295 9276 19329 9676
rect 19329 9276 19338 9676
rect 19128 7700 19137 8100
rect 19137 7700 19171 8100
rect 19171 7700 19180 8100
rect 19602 9276 19611 9676
rect 19611 9276 19645 9676
rect 19645 9276 19654 9676
rect 19444 7700 19453 8100
rect 19453 7700 19487 8100
rect 19487 7700 19496 8100
rect 19918 9276 19927 9676
rect 19927 9276 19961 9676
rect 19961 9276 19970 9676
rect 19760 7700 19769 8100
rect 19769 7700 19803 8100
rect 19803 7700 19812 8100
rect 20291 9737 20400 9935
rect 20400 9737 20413 10277
rect 20076 7700 20085 8100
rect 20085 7700 20119 8100
rect 20119 7700 20128 8100
rect 20261 7473 20274 9488
rect 20274 7473 20383 9488
rect 20261 7444 20383 7473
rect 18343 7373 20383 7444
rect 18343 7290 20384 7373
rect 18343 7243 20160 7290
rect 16178 7180 16230 7183
rect 16178 6783 16185 7180
rect 16185 6783 16223 7180
rect 16223 6783 16230 7180
rect 16693 7177 16869 7186
rect 16693 7143 16869 7177
rect 16693 7134 16869 7143
rect 17279 7177 17455 7186
rect 17279 7143 17455 7177
rect 17279 7134 17455 7143
rect 17865 7177 18041 7186
rect 17865 7143 18041 7177
rect 17865 7134 18041 7143
rect 16169 6521 16239 6539
rect 16169 6124 16185 6521
rect 16185 6124 16223 6521
rect 16223 6124 16239 6521
rect 16169 6107 16239 6124
rect 18519 6378 19526 6561
rect 18082 5147 18091 5657
rect 18091 5147 18125 5657
rect 18125 5147 18134 5657
rect 16693 5119 16869 5128
rect 16693 5085 16869 5119
rect 16693 5076 16869 5085
rect 17279 5119 17455 5128
rect 17279 5085 17455 5119
rect 17279 5076 17455 5085
rect 17865 5119 18041 5128
rect 17865 5085 18041 5119
rect 17865 5076 18041 5085
rect 16693 4715 16869 4724
rect 16693 4681 16869 4715
rect 16693 4672 16869 4681
rect 17279 4715 17455 4724
rect 17279 4681 17455 4715
rect 17279 4672 17455 4681
rect 17865 4715 18041 4724
rect 17865 4681 18041 4715
rect 17865 4672 18041 4681
rect 18082 2685 18091 3185
rect 18091 2685 18125 3185
rect 18125 2685 18134 3185
rect 16693 2657 16869 2666
rect 16693 2623 16869 2657
rect 16693 2614 16869 2623
rect 17279 2657 17455 2666
rect 17279 2623 17455 2657
rect 17279 2614 17455 2623
rect 17865 2657 18041 2666
rect 17865 2623 18041 2657
rect 17865 2614 18041 2623
rect 18714 3022 18784 3039
rect 18714 2625 18730 3022
rect 18730 2625 18768 3022
rect 18768 2625 18784 3022
rect 18714 2607 18784 2625
rect 19602 3022 19673 3039
rect 19602 2625 19618 3022
rect 19618 2625 19656 3022
rect 19656 2625 19673 3022
rect 19602 2607 19673 2625
rect 20099 2391 20160 7243
rect 20160 2391 20384 7290
rect 13755 2263 16522 2384
rect 16918 2263 18007 2384
rect 18209 2263 18322 2384
rect 20099 2380 20384 2391
rect 18651 2259 20384 2380
rect 21320 8161 24092 8164
rect 21320 8145 21325 8161
rect 21325 8145 24025 8161
rect 21195 8129 24025 8145
rect 24025 8129 24092 8161
rect 21195 8031 24090 8129
rect 21195 3591 21504 8031
rect 21504 8022 23911 8031
rect 23911 8022 24090 8031
rect 24090 8022 24092 8129
rect 23005 7945 23725 7954
rect 23005 7911 23725 7945
rect 23005 7902 23725 7911
rect 21654 6127 21665 7127
rect 21665 6127 21699 7127
rect 21699 6127 21710 7127
rect 24395 8159 25879 8168
rect 24395 8149 26789 8159
rect 26789 8149 26835 8159
rect 24395 8040 26835 8149
rect 21749 6087 22469 6096
rect 21749 6053 22469 6087
rect 21749 6044 22469 6053
rect 21979 5795 23721 5958
rect 21749 5695 22469 5704
rect 21749 5661 22469 5695
rect 21749 5652 22469 5661
rect 21654 5285 21665 5608
rect 21665 5285 21699 5608
rect 21699 5285 21710 5608
rect 21653 3865 21665 4865
rect 21665 3865 21699 4865
rect 21699 3865 21709 4865
rect 23909 4060 23911 7809
rect 23911 4311 24090 7809
rect 24090 4311 24092 7809
rect 24843 7945 25413 7954
rect 24843 7911 25413 7945
rect 24843 7902 25413 7911
rect 24364 5025 24618 7772
rect 25049 7687 25619 7696
rect 25049 7653 25619 7687
rect 25049 7644 25619 7653
rect 25836 7537 26835 8040
rect 24883 7369 26835 7537
rect 24883 7354 25918 7369
rect 24843 7239 25563 7248
rect 24843 7205 25563 7239
rect 24843 7196 25563 7205
rect 25799 6981 26519 6990
rect 25799 6947 26519 6981
rect 25799 6938 26519 6947
rect 24843 6723 25563 6732
rect 24843 6689 25563 6723
rect 24843 6680 25563 6689
rect 25799 6465 26519 6474
rect 25799 6431 26519 6465
rect 25799 6422 26519 6431
rect 24843 6207 25563 6216
rect 24843 6173 25563 6207
rect 24843 6164 25563 6173
rect 25799 5949 26519 5958
rect 25799 5915 26519 5949
rect 25799 5906 26519 5915
rect 24843 5691 25563 5700
rect 24843 5657 25563 5691
rect 24843 5648 25563 5657
rect 26708 5601 26835 7369
rect 25800 5433 26520 5442
rect 25800 5399 26519 5433
rect 26519 5399 26520 5433
rect 25800 5390 26520 5399
rect 24739 5203 24750 5371
rect 24750 5203 24784 5371
rect 24784 5203 24795 5371
rect 24843 5175 25563 5184
rect 24843 5141 25563 5175
rect 24843 5132 25563 5141
rect 26709 5025 26835 5334
rect 24358 4469 26835 5025
rect 26835 4492 26836 5334
rect 23911 4060 26905 4311
rect 23909 4053 24020 4060
rect 24020 4050 26905 4060
rect 23005 3837 23725 3846
rect 23005 3803 23725 3837
rect 23005 3794 23725 3803
rect 24678 3837 25398 3846
rect 24678 3803 25398 3837
rect 24678 3794 25398 3803
rect 21195 3233 24301 3591
rect 21199 3201 24301 3233
rect 21199 3147 24290 3201
rect 24290 3147 24295 3201
rect 21199 3106 24295 3147
rect 21437 2715 21446 2915
rect 21446 2715 21480 2915
rect 21480 2715 21489 2915
rect 21023 2035 21199 2403
rect 21199 2035 21328 2403
rect 21695 1939 21704 2139
rect 21704 1939 21738 2139
rect 21738 1939 21747 2139
rect 21508 1889 21639 1898
rect 21953 2715 21962 2915
rect 21962 2715 21996 2915
rect 21996 2715 22005 2915
rect 22211 1939 22220 2139
rect 22220 1939 22254 2139
rect 22254 1939 22263 2139
rect 22469 2715 22478 2915
rect 22478 2715 22512 2915
rect 22512 2715 22521 2915
rect 22727 1939 22736 2139
rect 22736 1939 22770 2139
rect 22770 1939 22779 2139
rect 22985 2715 22994 2915
rect 22994 2715 23028 2915
rect 23028 2715 23037 2915
rect 23243 1939 23252 2139
rect 23252 1939 23286 2139
rect 23286 1939 23295 2139
rect 23501 2715 23510 2915
rect 23510 2715 23544 2915
rect 23544 2715 23553 2915
rect 23759 1939 23768 2139
rect 23768 1939 23802 2139
rect 23802 1939 23811 2139
rect 24017 2715 24026 2915
rect 24026 2715 24060 2915
rect 24060 2715 24069 2915
rect 21508 1855 21639 1889
rect 21508 1846 21639 1855
rect 24187 2035 24295 3106
rect 24187 1784 24295 1868
rect 24578 2815 24594 3715
rect 24594 2815 24628 3715
rect 24628 2815 24642 3715
rect 24678 1979 25398 1987
rect 24678 1945 25398 1979
rect 24678 1935 25398 1945
rect 26479 1854 26830 1855
rect 26830 1854 26905 4050
rect 21215 1656 24295 1784
rect 24549 1663 26899 1854
rect 26899 1663 26905 1854
<< metal2 >>
rect 2433 42578 5829 42588
rect 2046 30457 2433 30467
rect 2688 42337 5603 42347
rect 5815 42337 5829 42347
rect 6032 31303 10883 31313
rect 6032 31108 10759 31118
rect 5603 30990 5815 31000
rect 10602 30906 10666 30916
rect 6224 30830 6276 30840
rect 2784 30766 2856 30776
rect 2784 30356 2856 30366
rect 5459 30763 6224 30773
rect 5511 30730 6224 30763
rect 10602 30796 10666 30806
rect 5511 30713 6276 30730
rect 6295 30679 6548 30689
rect 6295 30612 6548 30622
rect 10229 30686 10589 30696
rect 10229 30603 10589 30613
rect 5459 30356 5511 30366
rect 6031 30536 10759 30546
rect 10874 31108 10883 31118
rect 10874 30536 10882 30546
rect 10882 30351 10889 30408
rect 6031 30341 10889 30351
rect 2688 30250 5815 30260
rect 2446 30057 5815 30063
rect 2046 30053 5815 30057
rect 10489 30171 10889 30341
rect 25088 30171 25439 30181
rect 2046 30047 2446 30053
rect 10489 29859 25088 30171
rect 25088 29849 25439 29859
rect 11068 29793 11226 29803
rect 11068 29294 11226 29599
rect 4796 29136 11226 29294
rect 4796 14947 4954 29136
rect 6236 27983 7095 27993
rect 13986 27818 14066 27828
rect 12861 27808 13986 27818
rect 13258 27756 13986 27808
rect 12861 27746 13986 27756
rect 6236 27572 7095 27582
rect 13986 27334 14066 27344
rect 15378 26070 15907 26080
rect 15378 25974 15907 25984
rect 12958 25144 13258 25154
rect 12958 25082 13258 25092
rect 5742 24624 5981 24631
rect 5742 24621 11232 24624
rect 5981 24614 11232 24621
rect 11232 24599 12844 24609
rect 11232 24198 12844 24204
rect 5981 24194 12844 24198
rect 5981 24188 11232 24194
rect 7152 24120 8168 24130
rect 6180 24112 6240 24120
rect 6180 24110 6710 24112
rect 6240 24102 6710 24110
rect 6240 24068 6650 24102
rect 6180 24040 6240 24050
rect 7212 24068 7638 24120
rect 7698 24068 8108 24120
rect 7152 24058 7212 24068
rect 7638 24058 7698 24068
rect 8108 24058 8168 24068
rect 8610 24120 9140 24130
rect 8670 24068 9080 24120
rect 8610 24058 8670 24068
rect 9080 24058 9140 24068
rect 9582 24120 10112 24130
rect 9642 24068 10052 24120
rect 9582 24058 9642 24068
rect 10052 24058 10112 24068
rect 10554 24120 10614 24188
rect 10554 24058 10614 24068
rect 6650 24040 6710 24050
rect 6280 23961 6332 23971
rect 6558 23961 6610 23971
rect 6332 23860 6558 23961
rect 6280 22951 6332 22961
rect 6558 22951 6610 22961
rect 6768 23963 6820 23971
rect 7046 23963 7098 23973
rect 6768 23961 7046 23963
rect 6820 23862 7046 23961
rect 6768 22951 6820 22961
rect 7046 22953 7098 22963
rect 7737 23966 7789 23976
rect 8016 23966 8068 23976
rect 7789 23865 8016 23966
rect 7737 22956 7789 22966
rect 8016 22956 8068 22966
rect 8225 23964 8277 23974
rect 8500 23964 8552 23974
rect 8277 23863 8500 23964
rect 8225 22954 8277 22964
rect 8500 22954 8552 22964
rect 8712 23963 8764 23973
rect 8987 23963 9039 23973
rect 8764 23862 8987 23963
rect 8712 22953 8764 22963
rect 8987 22953 9039 22963
rect 9197 23964 9249 23973
rect 9473 23964 9525 23973
rect 9197 23963 9525 23964
rect 9684 23963 9736 23973
rect 9959 23963 10011 23973
rect 9249 23863 9473 23963
rect 9197 22953 9249 22963
rect 9682 23862 9684 23963
rect 9473 22953 9525 22963
rect 9736 23862 9959 23963
rect 9684 22953 9736 22963
rect 9959 22953 10011 22963
rect 10169 23972 10221 23973
rect 10446 23972 10498 23973
rect 10169 23963 10498 23972
rect 10221 23871 10446 23963
rect 10169 22953 10221 22963
rect 13158 23617 13258 25082
rect 15564 24057 20117 24059
rect 15564 24049 20149 24057
rect 20117 24047 20149 24049
rect 15564 23788 19697 23789
rect 15564 23779 20149 23788
rect 19697 23778 20149 23779
rect 10446 22953 10498 22963
rect 10823 23607 15840 23617
rect 10823 23517 15788 23607
rect 10823 21049 10903 23517
rect 15788 23397 15840 23407
rect 19846 23607 19898 23617
rect 19898 23407 20433 23497
rect 19846 23397 20433 23407
rect 11332 22831 11384 22841
rect 11055 22631 11332 22721
rect 11055 22621 11384 22631
rect 15388 22831 15444 22841
rect 15444 22631 20211 22721
rect 15388 22621 20211 22631
rect 11055 21955 11155 22621
rect 16147 22381 20041 22391
rect 11352 22356 15126 22366
rect 11352 22162 15126 22172
rect 16147 22136 20041 22146
rect 11055 21945 11209 21955
rect 20111 21945 20211 22621
rect 11055 21845 11109 21945
rect 11209 21935 15840 21945
rect 11209 21845 15788 21935
rect 11109 21835 11209 21845
rect 11339 21159 11391 21169
rect 10823 20959 11339 21049
rect 10823 20949 11391 20959
rect 11279 20783 15029 20793
rect 11279 20686 15029 20696
rect 15105 20291 15181 21845
rect 15530 21768 15686 21778
rect 15788 21725 15840 21735
rect 19846 21935 20211 21945
rect 19898 21845 20211 21935
rect 19846 21725 19898 21735
rect 19961 21752 20148 21762
rect 15686 21187 19961 21197
rect 15397 21159 15449 21169
rect 15530 21151 15537 21161
rect 15537 21100 20148 21110
rect 20127 21049 20227 21059
rect 20333 21049 20433 23397
rect 15449 20959 20127 21049
rect 15397 20949 20127 20959
rect 20227 20949 20433 21049
rect 20127 20939 20227 20949
rect 15105 20215 20987 20291
rect 5742 19767 5981 19777
rect 6180 20050 6240 20060
rect 6180 19697 6240 19998
rect 6666 20044 6726 20054
rect 7136 20044 7196 20054
rect 6726 19992 7136 20044
rect 6666 19982 7196 19992
rect 7622 20044 7682 20054
rect 6169 19687 6246 19697
rect 6169 19577 6246 19587
rect 5273 19462 5373 19472
rect 7622 19462 7682 19992
rect 8124 20044 8184 20054
rect 8594 20044 8654 20054
rect 8184 19992 8594 20044
rect 8124 19982 8654 19992
rect 9096 20044 9156 20054
rect 9566 20044 9626 20054
rect 9156 19992 9566 20044
rect 9096 19982 9626 19992
rect 10068 20044 10128 20054
rect 10538 20044 10598 20054
rect 10128 19992 10538 20044
rect 10068 19982 10598 19992
rect 5373 19410 7682 19462
rect 5273 19375 5373 19385
rect 6349 19039 6401 19410
rect 9350 19143 10350 19153
rect 9350 19077 10350 19087
rect 11506 19143 12506 19153
rect 11506 19077 12506 19087
rect 6349 18503 6401 18763
rect 6349 18217 6401 18227
rect 10407 19039 10459 19049
rect 10407 18503 10459 18763
rect 19815 19039 19879 19049
rect 20911 18780 20987 20215
rect 20911 18718 20987 18728
rect 21403 18796 21503 18806
rect 21403 18722 21503 18732
rect 19815 18429 19879 18439
rect 21035 18700 21091 18710
rect 6342 17639 6406 17649
rect 6342 17429 6406 17439
rect 10407 17639 10459 18227
rect 21035 17690 21091 17700
rect 21539 18658 21595 18668
rect 4796 14937 9420 14947
rect 4796 14885 8420 14937
rect 4796 14875 9420 14885
rect 4796 12094 4954 14875
rect 10407 14835 10459 17063
rect 11431 17663 11495 17673
rect 21539 17648 21595 17658
rect 11431 17053 11495 17063
rect 15495 17563 15547 17573
rect 11431 16635 11495 16645
rect 15495 16635 15547 17063
rect 15495 16125 15547 16135
rect 15763 17563 15815 17573
rect 15763 16635 15815 17063
rect 15763 16125 15815 16135
rect 11431 16025 11495 16035
rect 19815 15259 19879 15269
rect 8054 14789 8246 14799
rect 8349 14786 8401 14796
rect 8246 14659 8349 14729
rect 8246 14649 8401 14659
rect 15495 14850 15547 14860
rect 10459 14659 15495 14733
rect 15763 14850 15815 14860
rect 15547 14659 15763 14733
rect 19805 14792 19815 14810
rect 19879 14792 19889 14810
rect 19805 14778 19889 14792
rect 15815 14716 21530 14733
rect 15815 14664 20911 14716
rect 20987 14664 21415 14716
rect 21491 14664 21530 14716
rect 15815 14659 21530 14664
rect 10407 14649 21530 14659
rect 21526 14480 22053 14481
rect 21513 14474 22053 14480
rect 8246 14471 22054 14474
rect 8246 14464 21526 14471
rect 22053 14464 22054 14471
rect 8054 14440 8056 14450
rect 7961 14001 8056 14232
rect 7961 13991 21526 14001
rect 21513 13979 21526 13991
rect 22053 13979 22054 13980
rect 21526 13970 22054 13979
rect 21526 13969 22053 13970
rect 9591 13059 10125 13069
rect 9591 12834 10125 12927
rect 7800 12824 10813 12834
rect 10778 12724 10813 12824
rect 10778 12663 10779 12673
rect 7800 12509 10284 12519
rect 8064 12335 8116 12509
rect 8064 12125 8116 12135
rect 10122 12311 10174 12321
rect 4796 12084 8844 12094
rect 4796 12032 8135 12084
rect 4796 12022 8844 12032
rect 5836 11969 10075 11979
rect 5983 11751 10075 11761
rect 5836 11184 5983 11194
rect 6051 11548 6122 11558
rect 10122 11548 10174 12135
rect 6051 11162 6122 11172
rect 9770 11172 10122 11214
rect 9770 11162 10174 11172
rect 5273 11125 5373 11135
rect 5373 11115 7135 11125
rect 5373 11063 6135 11115
rect 5373 11053 7135 11063
rect 5273 11043 5373 11053
rect 5840 10956 9712 10966
rect 5840 10830 7787 10840
rect 6170 10562 6234 10572
rect 6170 10316 6234 10326
rect 7644 10322 7708 10332
rect 6892 10194 6985 10204
rect 7644 10076 7708 10086
rect 6892 9960 6985 9970
rect 4365 9919 4498 9929
rect 4498 9918 5684 9919
rect 6235 9918 6335 9928
rect 7171 9918 7271 9928
rect 4498 9818 6235 9918
rect 6335 9818 7171 9918
rect 4365 9808 4498 9818
rect 6235 9808 6335 9818
rect 7171 9808 7271 9818
rect 3925 9768 4058 9778
rect 6607 9768 6707 9778
rect 7549 9768 7649 9778
rect 4058 9668 6607 9768
rect 6707 9668 7549 9768
rect 3925 9658 4058 9668
rect 6607 9658 6707 9668
rect 7549 9658 7649 9668
rect 7644 9520 7708 9530
rect 6170 9280 6234 9290
rect 7644 9275 7708 9285
rect 6170 9034 6234 9044
rect 5870 8871 7787 8881
rect 7942 10830 8812 10840
rect 7942 8871 7960 8881
rect 5870 8757 7960 8767
rect 8950 10830 9712 10840
rect 9770 10782 9836 11162
rect 12349 12101 12894 12111
rect 12349 11127 12894 11926
rect 13324 11262 20778 11398
rect 11880 11124 13004 11127
rect 10284 10796 10655 10806
rect 9580 10730 10026 10782
rect 9580 10580 9632 10730
rect 9036 10304 9100 10314
rect 9036 10094 9100 10104
rect 9036 9495 9100 9505
rect 9036 9285 9100 9295
rect 9580 9495 9632 10380
rect 9580 9285 9632 9295
rect 9974 10580 10026 10730
rect 9974 9495 10026 10380
rect 10506 10580 10570 10590
rect 10506 10370 10570 10380
rect 9974 9285 10026 9295
rect 10506 9219 10570 9229
rect 10506 9009 10570 9019
rect 8950 8863 10655 8873
rect 10776 10796 10779 10806
rect 11848 11117 13004 11124
rect 11848 11114 11880 11117
rect 12899 11079 13004 11117
rect 11967 10996 12773 11006
rect 12340 10853 12392 10996
rect 11848 10394 11967 10404
rect 12024 10777 12076 10787
rect 12340 10743 12392 10753
rect 12656 10777 12708 10787
rect 11366 10242 11466 10252
rect 12024 10226 12076 10677
rect 12131 10349 12206 10355
rect 12656 10349 12708 10677
rect 12901 10996 13004 11079
rect 12773 10408 12901 10418
rect 13324 10349 13473 11262
rect 20291 11042 20413 11050
rect 12131 10295 12148 10349
rect 12203 10295 13473 10349
rect 12131 10289 12206 10295
rect 12321 10226 12394 10232
rect 11466 10172 12330 10226
rect 12384 10172 12394 10226
rect 11366 10162 11466 10172
rect 11241 9898 11310 9908
rect 12122 9649 12174 10172
rect 12321 10166 12394 10172
rect 11447 9648 12174 9649
rect 11408 9638 12174 9648
rect 11460 9597 12122 9638
rect 11408 9548 11460 9558
rect 11566 9542 11618 9552
rect 11964 9542 12016 9552
rect 12122 9548 12174 9558
rect 12520 9648 12572 10295
rect 13324 10293 13473 10295
rect 13755 11040 20413 11042
rect 13755 11032 20291 11040
rect 13384 9900 13448 9910
rect 12520 9638 13286 9648
rect 12572 9596 13234 9638
rect 12520 9548 12572 9558
rect 11618 9462 11964 9508
rect 11566 9297 11618 9462
rect 11964 9452 12016 9462
rect 12678 9542 12730 9552
rect 13076 9542 13128 9552
rect 13234 9548 13286 9558
rect 12730 9462 13076 9498
rect 12678 9452 13128 9462
rect 12035 9412 12103 9422
rect 12035 9346 12103 9356
rect 12678 9297 12730 9452
rect 13147 9412 13215 9422
rect 13147 9346 13215 9356
rect 11310 9287 13384 9297
rect 11230 9173 11241 9271
rect 13446 9277 13448 9287
rect 11230 9163 13446 9173
rect 8812 8737 8821 8741
rect 8812 8731 10655 8737
rect 8821 8728 10655 8731
rect 8821 8727 10776 8728
rect 10655 8718 10776 8727
rect 8523 8650 8589 8660
rect 5318 8640 8523 8650
rect 5295 8630 5318 8640
rect 8589 8626 10790 8636
rect 11237 8566 11709 9163
rect 4528 8529 4703 8539
rect 4703 8129 5295 8529
rect 4528 8119 4703 8129
rect 5375 8550 8523 8560
rect 5450 8387 5514 8397
rect 5450 8313 5514 8323
rect 6714 8387 6766 8550
rect 6714 8277 6766 8287
rect 7112 8387 7164 8550
rect 7112 8277 7164 8287
rect 8364 8275 8428 8285
rect 8364 8201 8428 8211
rect 5375 8009 8523 8019
rect 8589 8554 8824 8564
rect 8589 7995 8824 8005
rect 8961 8554 9704 8564
rect 9036 8387 9100 8397
rect 9036 8277 9100 8287
rect 9540 8311 9592 8321
rect 9113 8171 9273 8181
rect 9113 8097 9273 8107
rect 9540 8005 9592 8211
rect 8961 7995 9704 8005
rect 9897 8554 10665 8564
rect 10014 8388 10066 8554
rect 10014 8278 10066 8288
rect 10506 8388 10570 8398
rect 10506 8278 10570 8288
rect 10085 8173 10245 8183
rect 10085 8099 10245 8109
rect 9897 7995 10665 8005
rect 10790 8094 11709 8566
rect 10790 7995 10802 8005
rect 8589 7923 10802 7933
rect 5375 7859 8523 7869
rect 5450 7671 5514 7681
rect 5450 7597 5514 7607
rect 6714 7595 6766 7605
rect 6714 7305 6766 7495
rect 7112 7595 7164 7605
rect 7112 7305 7164 7495
rect 8364 7548 8428 7558
rect 8364 7474 8428 7484
rect 5375 7295 8523 7305
rect 5375 7145 8523 7155
rect 5450 6955 5514 6965
rect 5450 6881 5514 6891
rect 8364 6955 8428 6965
rect 6714 6879 6766 6889
rect 6714 6574 6766 6779
rect 7112 6879 7164 6889
rect 8364 6881 8428 6891
rect 7112 6574 7164 6779
rect 5375 6564 8523 6574
rect 5375 6414 8523 6424
rect 8364 6239 8428 6249
rect 6714 6163 6766 6173
rect 5450 6127 5514 6137
rect 5450 6053 5514 6063
rect 6714 5877 6766 6063
rect 7112 6163 7164 6173
rect 8364 6165 8428 6175
rect 7112 5877 7164 6063
rect 5375 5867 8523 5877
rect 5272 5730 5295 5825
rect 5272 5727 5335 5730
rect 5272 5720 8523 5727
rect 5272 5717 8589 5720
rect 8523 5710 8589 5717
rect 13750 2396 13755 2406
rect 13869 10854 16576 10864
rect 16576 9925 20291 9935
rect 20291 9727 20413 9737
rect 18022 9686 18074 9687
rect 20642 9686 20778 11262
rect 16133 9677 20778 9686
rect 16133 9676 18022 9677
rect 16133 9550 16758 9676
rect 16133 7183 16274 9550
rect 16810 9550 17074 9676
rect 16758 9266 16810 9276
rect 17126 9550 17390 9676
rect 17074 9266 17126 9276
rect 17442 9550 17706 9676
rect 17390 9266 17442 9276
rect 17758 9550 18022 9676
rect 17706 9266 17758 9276
rect 18074 9676 20778 9677
rect 18074 9550 18338 9676
rect 18022 9267 18074 9277
rect 18390 9550 18654 9676
rect 18338 9266 18390 9276
rect 18706 9550 18970 9676
rect 18654 9266 18706 9276
rect 19022 9550 19286 9676
rect 18970 9266 19022 9276
rect 19338 9550 19602 9676
rect 19286 9266 19338 9276
rect 19654 9550 19918 9676
rect 19602 9266 19654 9276
rect 19970 9550 20778 9676
rect 19918 9266 19970 9276
rect 20261 9488 20383 9498
rect 16133 6783 16178 7183
rect 16230 6783 16274 7183
rect 16600 8100 16652 8110
rect 16916 8100 16968 8110
rect 16652 7700 16916 7826
rect 17232 8100 17284 8110
rect 16968 7700 17232 7826
rect 17548 8100 17600 8110
rect 17284 7700 17548 7826
rect 17864 8100 17916 8110
rect 17600 7700 17864 7826
rect 18180 8100 18232 8110
rect 17916 7700 18180 7826
rect 18496 8100 18548 8110
rect 18232 7700 18496 7826
rect 18812 8100 18864 8110
rect 18548 7700 18812 7826
rect 19128 8100 19180 8110
rect 18864 7700 19128 7826
rect 19444 8100 19496 8110
rect 19180 7700 19444 7826
rect 19760 8100 19812 8110
rect 19496 7700 19760 7826
rect 20076 8100 20128 8110
rect 19812 7700 20076 7826
rect 16600 7690 20128 7700
rect 16600 7196 16652 7690
rect 18343 7444 20261 7454
rect 21320 8164 24092 8174
rect 21195 8145 21320 8155
rect 24395 8169 25879 8178
rect 26466 8169 26867 8178
rect 24395 8168 26933 8169
rect 25879 8159 26466 8168
rect 24395 8030 25836 8040
rect 20383 7373 20384 7383
rect 18343 7233 20099 7243
rect 16600 7186 16881 7196
rect 16600 7134 16693 7186
rect 16869 7134 16881 7186
rect 16600 7124 16881 7134
rect 17267 7186 18041 7196
rect 17267 7134 17279 7186
rect 17455 7134 17865 7186
rect 17267 7124 18041 7134
rect 16133 6773 16274 6783
rect 18519 6561 20099 6571
rect 16169 6539 16239 6549
rect 16168 6107 16169 6200
rect 19526 6378 20099 6561
rect 18519 6368 20099 6378
rect 19496 6367 20099 6368
rect 16239 6107 16240 6200
rect 16168 4734 16240 6107
rect 18082 5657 18134 5667
rect 18134 5147 18460 5193
rect 18082 5141 18460 5147
rect 17865 5138 18041 5141
rect 16693 5128 17475 5138
rect 16869 5076 17279 5128
rect 17455 5076 17475 5128
rect 16693 5066 17475 5076
rect 17853 5131 18045 5138
rect 17853 5073 17865 5131
rect 18041 5073 18045 5131
rect 17853 5066 18045 5073
rect 17865 5063 18041 5066
rect 16168 4724 16888 4734
rect 16168 4672 16693 4724
rect 16869 4672 16888 4724
rect 16168 4662 16888 4672
rect 17259 4724 18041 4734
rect 17259 4672 17279 4724
rect 17455 4672 17865 4724
rect 17259 4662 18041 4672
rect 18082 3185 18134 3195
rect 17865 2676 18041 2679
rect 16693 2666 17471 2676
rect 16869 2614 17279 2666
rect 17455 2614 17471 2666
rect 16693 2604 17471 2614
rect 17853 2669 18041 2676
rect 17853 2611 17865 2669
rect 17853 2604 18041 2611
rect 17865 2601 18041 2604
rect 13869 2396 16043 2406
rect 13607 2253 13750 2394
rect 16043 2384 16546 2394
rect 16522 2263 16546 2384
rect 16043 2253 16546 2263
rect 16896 2384 18007 2394
rect 16896 2263 16918 2384
rect 16896 2253 18007 2263
rect 13750 2171 16043 2181
rect 11778 678 11958 688
rect 18082 678 18134 2685
rect 18209 2384 18322 2394
rect 18209 2253 18322 2263
rect 11768 626 11778 678
rect 11958 626 18134 678
rect 11778 601 11958 611
rect 15642 455 15822 465
rect 18408 455 18460 5141
rect 18714 3039 18784 3049
rect 18714 2597 18784 2607
rect 19602 3039 19673 3049
rect 19602 2597 19673 2607
rect 18624 2380 20099 2390
rect 21504 8012 24092 8022
rect 23005 7954 25413 7964
rect 23725 7902 24843 7954
rect 23005 7892 25413 7902
rect 23909 7809 24092 7819
rect 21654 7127 21710 7137
rect 21654 5608 21710 6127
rect 21749 6096 22469 6106
rect 21749 6034 22469 6044
rect 21749 5714 21917 6034
rect 21979 5962 23721 5968
rect 21979 5958 23909 5962
rect 23721 5795 23909 5958
rect 21979 5785 23721 5795
rect 21749 5704 22469 5714
rect 21749 5642 22469 5652
rect 21654 4875 21710 5285
rect 21653 4865 21710 4875
rect 21709 4862 21710 4865
rect 24364 7772 24618 7782
rect 24358 5025 24364 5035
rect 25049 7696 25619 7706
rect 25049 7634 25619 7644
rect 25410 7547 25619 7634
rect 26867 8078 26933 8168
rect 24618 7537 25836 7547
rect 26835 7607 26867 7617
rect 24618 7354 24883 7537
rect 25918 7359 26708 7369
rect 24618 7344 25918 7354
rect 25352 7258 25563 7344
rect 24843 7248 25563 7258
rect 24843 7186 25563 7196
rect 24843 6742 24990 7186
rect 25799 6990 26519 7000
rect 26519 6938 26520 6972
rect 25799 6928 26520 6938
rect 24843 6732 25563 6742
rect 24843 6670 25563 6680
rect 24843 6226 24990 6670
rect 26348 6484 26520 6928
rect 25799 6474 26520 6484
rect 26519 6422 26520 6474
rect 25799 6412 26520 6422
rect 24843 6216 25563 6226
rect 24843 6154 25563 6164
rect 24843 5710 24990 6154
rect 26348 5968 26520 6412
rect 25799 5958 26520 5968
rect 26519 5906 26520 5958
rect 25799 5896 26520 5906
rect 24843 5700 25563 5710
rect 24843 5638 25563 5648
rect 24739 5371 24795 5381
rect 24739 5193 24795 5203
rect 24843 5194 24990 5638
rect 26348 5535 26520 5896
rect 26708 5591 26835 5601
rect 27234 5535 27414 5545
rect 26348 5452 27234 5535
rect 25800 5442 27234 5452
rect 26520 5390 27234 5442
rect 25800 5380 27234 5390
rect 27234 5370 27414 5380
rect 26709 5334 26836 5344
rect 24843 5184 25563 5194
rect 24843 5122 25563 5132
rect 24843 5035 24990 5122
rect 24618 5025 26709 5035
rect 26835 4482 26836 4492
rect 24358 4459 26835 4469
rect 24092 4311 26905 4321
rect 23909 4050 24020 4053
rect 23909 4043 26830 4050
rect 24020 4040 26830 4043
rect 21653 3855 21709 3865
rect 23005 3846 25398 3856
rect 23725 3794 24678 3846
rect 23005 3784 25398 3794
rect 24578 3715 24642 3725
rect 21504 3591 24301 3601
rect 21113 3259 21167 3260
rect 21113 3233 21195 3259
rect 21113 3106 21199 3233
rect 24295 3191 24301 3201
rect 21113 3096 24187 3106
rect 21437 2925 21513 3096
rect 21954 2925 22046 3096
rect 22438 2925 22530 3096
rect 22980 2925 23071 3096
rect 23494 2925 23585 3096
rect 24011 2925 24102 3096
rect 21437 2915 24102 2925
rect 21489 2873 21953 2915
rect 21437 2705 21489 2715
rect 22005 2873 22469 2915
rect 21953 2705 22005 2715
rect 22521 2873 22985 2915
rect 22469 2705 22521 2715
rect 23037 2873 23501 2915
rect 22985 2705 23037 2715
rect 23553 2873 24017 2915
rect 23501 2705 23553 2715
rect 24069 2914 24102 2915
rect 24017 2705 24069 2715
rect 18624 2259 18651 2380
rect 18624 2249 20384 2259
rect 21023 2403 21328 2413
rect 18704 2087 18794 2097
rect 21023 2025 21328 2035
rect 21695 2139 21747 2149
rect 18704 1908 18794 1988
rect 22211 2139 22263 2149
rect 21747 1939 22211 1998
rect 22727 2139 22779 2149
rect 22263 1939 22727 1998
rect 23243 2139 23295 2149
rect 22779 1939 23243 1998
rect 23759 2139 23811 2149
rect 23295 1939 23759 1998
rect 24578 2805 24642 2815
rect 24187 2027 24295 2035
rect 23811 1987 25403 1998
rect 23811 1939 24678 1987
rect 21695 1935 24678 1939
rect 25398 1935 25403 1987
rect 21695 1926 25403 1935
rect 18704 1898 21639 1908
rect 18704 1846 21508 1898
rect 18704 1836 21639 1846
rect 24187 1868 24295 1874
rect 19506 839 19687 1836
rect 21215 1784 24187 1794
rect 21215 1646 24295 1656
rect 24343 1577 24475 1926
rect 24678 1925 25398 1926
rect 26479 1864 26830 1865
rect 24549 1855 26830 1864
rect 24549 1854 26479 1855
rect 24549 1653 26905 1663
rect 24343 1418 24475 1428
rect 19506 680 19687 690
rect 15822 403 18460 455
rect 15642 385 15822 395
<< via2 >>
rect 2046 30250 2433 30457
rect 2433 30250 2446 30457
rect 2784 30366 2856 30766
rect 10602 30806 10666 30906
rect 6295 30622 6548 30679
rect 10229 30613 10589 30686
rect 2046 30063 2429 30250
rect 2429 30063 2446 30250
rect 5694 30156 5810 30233
rect 2046 30057 2446 30063
rect 25088 29859 25439 30171
rect 11068 29599 11226 29793
rect 6236 27582 7095 27983
rect 15378 25984 15907 26070
rect 6180 24102 6240 24110
rect 6180 24050 6240 24102
rect 19697 23789 20117 24047
rect 20117 23789 20149 24047
rect 19697 23788 20149 23789
rect 15388 22631 15390 22831
rect 15390 22631 15442 22831
rect 15442 22631 15444 22831
rect 11109 21845 11209 21945
rect 20127 20949 20227 21049
rect 6169 19587 6246 19687
rect 5273 19385 5373 19462
rect 9350 19087 10350 19143
rect 11506 19087 12506 19143
rect 19815 18439 19879 19039
rect 21403 18732 21503 18796
rect 6342 17439 6406 17639
rect 21035 17700 21091 18700
rect 11431 17063 11495 17663
rect 21539 17658 21595 18658
rect 11431 16035 11495 16635
rect 19815 14792 19879 15259
rect 21526 14464 22053 14471
rect 21526 14454 21806 14464
rect 21806 14454 22054 14464
rect 21526 14001 21822 14454
rect 21526 13991 21564 14001
rect 21564 13991 21822 14001
rect 21822 13991 22054 14454
rect 21526 13980 22054 13991
rect 21526 13979 22053 13980
rect 9591 12927 10125 13059
rect 6051 11172 6058 11548
rect 6058 11172 6116 11548
rect 6116 11172 6122 11548
rect 5273 11053 5373 11125
rect 6170 10327 6234 10562
rect 6170 10326 6234 10327
rect 6892 9970 6985 10194
rect 7644 10086 7708 10322
rect 4365 9818 4498 9919
rect 3925 9668 4058 9768
rect 6170 9044 6234 9280
rect 7644 9285 7708 9520
rect 12349 11926 12894 12101
rect 9036 10104 9100 10304
rect 9036 9295 9100 9495
rect 10506 10380 10570 10580
rect 10506 9019 10570 9219
rect 11366 10172 11466 10242
rect 12035 9356 12103 9412
rect 13147 9356 13215 9412
rect 4528 8129 4703 8529
rect 5450 8323 5514 8387
rect 8364 8211 8428 8275
rect 9036 8287 9100 8387
rect 9113 8107 9273 8171
rect 10506 8288 10570 8388
rect 10085 8109 10245 8173
rect 5450 7607 5514 7671
rect 8364 7484 8428 7548
rect 5450 6891 5514 6955
rect 8364 6891 8428 6955
rect 8364 6175 8428 6239
rect 5450 6063 5514 6127
rect 26466 8159 26867 8168
rect 17865 5128 18041 5131
rect 17865 5076 18041 5128
rect 17865 5073 18041 5076
rect 17865 2666 18041 2669
rect 17865 2614 18041 2666
rect 17865 2611 18041 2614
rect 13750 2263 13755 2396
rect 13755 2384 13869 2396
rect 13869 2384 16043 2396
rect 13755 2263 16043 2384
rect 13750 2181 16043 2263
rect 11778 611 11958 678
rect 18714 2607 18784 3039
rect 19602 2607 19673 3039
rect 21653 3865 21709 4865
rect 26466 7617 26835 8159
rect 26835 7617 26867 8159
rect 24739 5203 24795 5371
rect 27234 5380 27414 5535
rect 18704 1988 18794 2087
rect 21023 2035 21328 2403
rect 24578 2815 24642 3715
rect 24343 1428 24475 1577
rect 19506 690 19687 839
rect 15642 395 15822 455
<< metal3 >>
rect 11444 42754 17816 42782
rect 11444 36730 17732 42754
rect 17796 37227 17816 42754
rect 18340 42756 24712 42784
rect 18340 37227 24628 42756
rect 17796 36732 24628 37227
rect 24692 36732 24712 42756
rect 17796 36730 24712 36732
rect 11444 36704 24712 36730
rect 11444 36702 18680 36704
rect 17345 36326 18680 36702
rect 11443 36324 18680 36326
rect 11443 36298 24711 36324
rect 10592 30906 10693 30912
rect 10592 30806 10602 30906
rect 10666 30806 10693 30906
rect 10592 30801 10693 30806
rect 2774 30766 2866 30771
rect 2036 30457 2456 30462
rect 2036 30057 2046 30457
rect 2446 30057 2456 30457
rect 2774 30366 2784 30766
rect 2856 30366 2866 30766
rect 11443 30691 17731 36298
rect 10219 30686 17731 30691
rect 2774 30361 2866 30366
rect 6285 30679 6558 30684
rect 6285 30622 6295 30679
rect 6548 30622 6558 30679
rect 6285 30617 6558 30622
rect 2036 30052 2456 30057
rect 2784 29931 2856 30361
rect 5684 30233 5820 30238
rect 6285 30233 6364 30617
rect 10219 30613 10229 30686
rect 10589 30613 17731 30686
rect 10219 30608 17731 30613
rect 11443 30274 17731 30608
rect 17795 36296 24711 36298
rect 17795 35910 24627 36296
rect 17795 30274 17815 35910
rect 11443 30246 17815 30274
rect 18339 30272 24627 35910
rect 24691 30272 24711 36296
rect 18339 30244 24711 30272
rect 5684 30156 5694 30233
rect 5810 30156 6364 30233
rect 25078 30171 25449 30176
rect 5684 30151 5820 30156
rect 2769 13560 2869 29931
rect 25078 29859 25088 30171
rect 25439 29859 25449 30171
rect 25078 29854 25449 29859
rect 11058 29793 11236 29798
rect 11058 29599 11068 29793
rect 11226 29599 11236 29793
rect 11058 29594 11236 29599
rect 6226 27983 7105 27988
rect 6226 27582 6236 27983
rect 7095 27582 7105 27983
rect 6226 27577 7105 27582
rect 22064 27080 27936 27108
rect 15368 26070 15917 26075
rect 15368 25984 15378 26070
rect 15907 25984 15917 26070
rect 15368 25979 15917 25984
rect 5490 24045 5500 24115
rect 5598 24110 6250 24115
rect 5598 24050 6180 24110
rect 6240 24050 6250 24110
rect 5598 24045 6250 24050
rect 15378 22831 15454 25979
rect 19687 24050 20159 24052
rect 22064 24050 22084 27080
rect 19687 24047 22084 24050
rect 19687 23788 19697 24047
rect 20149 23790 22084 24047
rect 20149 23788 20159 23790
rect 19687 23783 20159 23788
rect 15378 22631 15388 22831
rect 15444 22631 15454 22831
rect 15378 22626 15454 22631
rect 11099 21945 11219 21950
rect 11099 21845 11109 21945
rect 11209 21845 11219 21945
rect 11099 21840 11219 21845
rect 22064 21556 22084 23790
rect 22148 21556 27936 27080
rect 22064 21528 27936 21556
rect 20117 21049 20237 21054
rect 20117 20949 20127 21049
rect 20227 20949 20237 21049
rect 20117 20944 20237 20949
rect 27101 20922 27832 21528
rect 22064 20894 27936 20922
rect 6159 19687 6256 19692
rect 6159 19587 6169 19687
rect 6246 19587 6256 19687
rect 6159 19582 6256 19587
rect 5263 19462 5383 19467
rect 5263 19385 5273 19462
rect 5373 19385 5383 19462
rect 5263 19380 5383 19385
rect 9340 19143 12516 19148
rect 9340 19087 9350 19143
rect 10350 19087 11506 19143
rect 12506 19087 12516 19143
rect 9340 19082 12516 19087
rect 19805 19039 19889 19044
rect 19805 18439 19815 19039
rect 19879 18439 19889 19039
rect 19805 18434 19889 18439
rect 21025 18796 21513 18808
rect 21025 18732 21403 18796
rect 21503 18732 21513 18796
rect 21025 18727 21513 18732
rect 21025 18726 21427 18727
rect 21025 18700 21101 18726
rect 21025 17700 21035 18700
rect 21091 17700 21101 18700
rect 22064 18663 22084 20894
rect 21025 17695 21101 17700
rect 21529 18658 22084 18663
rect 11421 17663 11505 17668
rect 6332 17639 6416 17644
rect 6332 17439 6342 17639
rect 6406 17439 6416 17639
rect 6332 17434 6416 17439
rect 11421 17063 11431 17663
rect 11495 17063 11505 17663
rect 21529 17658 21539 18658
rect 21595 18563 22084 18658
rect 21595 17658 21605 18563
rect 21529 17653 21605 17658
rect 11421 17058 11505 17063
rect 11421 16635 11505 16640
rect 11421 16035 11431 16635
rect 11495 16035 11505 16635
rect 11421 16030 11505 16035
rect 22064 15370 22084 18563
rect 22148 15370 27936 20894
rect 22064 15342 27936 15370
rect 19805 15259 19889 15264
rect 19805 14792 19815 15259
rect 19879 14792 19889 15259
rect 19805 14769 19889 14792
rect 21516 14471 22063 14476
rect 21516 13979 21526 14471
rect 22053 14469 22063 14471
rect 22053 14464 22064 14469
rect 22054 13980 22064 14464
rect 22053 13979 22064 13980
rect 21516 13975 22064 13979
rect 21516 13974 22063 13975
rect 2769 13460 11466 13560
rect 9581 13059 10135 13064
rect 9581 12927 9591 13059
rect 10125 12927 10135 13059
rect 9581 12922 10135 12927
rect 6041 11548 6132 11553
rect 6041 11172 6051 11548
rect 6122 11266 6132 11548
rect 6122 11172 6995 11266
rect 6041 11167 6995 11172
rect 6043 11166 6995 11167
rect 5263 11125 5383 11130
rect 5263 11053 5273 11125
rect 5373 11053 5383 11125
rect 5263 11048 5383 11053
rect 6160 10562 6244 10567
rect 6160 10326 6170 10562
rect 6234 10326 6244 10562
rect 6160 10321 6244 10326
rect 6882 10194 6995 11166
rect 8761 10580 10580 10585
rect 8761 10521 10506 10580
rect 6882 9970 6892 10194
rect 6985 9970 6995 10194
rect 7634 10322 7718 10327
rect 7634 10086 7644 10322
rect 7708 10181 7718 10322
rect 7708 10086 7981 10181
rect 7634 10081 7981 10086
rect 6882 9965 6995 9970
rect 4355 9919 4508 9924
rect 4355 9818 4365 9919
rect 4498 9818 4508 9919
rect 4355 9813 4508 9818
rect 3915 9768 4068 9773
rect 3915 9668 3925 9768
rect 4058 9668 4068 9768
rect 3915 9663 4068 9668
rect 7634 9520 7718 9525
rect 7634 9285 7644 9520
rect 7708 9285 7718 9520
rect 6160 9280 6244 9285
rect 7634 9280 7718 9285
rect 6160 9044 6170 9280
rect 6234 9139 6244 9280
rect 7881 9139 7981 10081
rect 8761 9500 8825 10521
rect 10496 10380 10506 10521
rect 10570 10380 10580 10580
rect 10496 10375 10580 10380
rect 9026 10304 9110 10309
rect 9026 10104 9036 10304
rect 9100 10104 9110 10304
rect 11366 10247 11466 13460
rect 12339 12101 12904 12106
rect 12339 11926 12349 12101
rect 12894 11926 12904 12101
rect 12339 11921 12904 11926
rect 11356 10242 11476 10247
rect 11356 10172 11366 10242
rect 11466 10172 11476 10242
rect 11356 10167 11476 10172
rect 9026 10099 9110 10104
rect 8761 9495 9110 9500
rect 8761 9436 9036 9495
rect 6234 9044 7981 9139
rect 6160 9039 7981 9044
rect 9026 9295 9036 9436
rect 9100 9295 9110 9495
rect 4518 8529 4713 8534
rect 2862 8129 2868 8529
rect 3266 8129 4528 8529
rect 4703 8129 4713 8529
rect 5439 8387 5587 8392
rect 6160 8388 6244 9039
rect 7633 8675 7643 8739
rect 7709 8675 7719 8739
rect 5439 8323 5450 8387
rect 5514 8323 5587 8387
rect 5439 8318 5587 8323
rect 6151 8322 6161 8388
rect 6244 8322 6254 8388
rect 7643 8255 7709 8675
rect 9026 8387 9110 9295
rect 12025 9412 12113 9417
rect 12025 9356 12035 9412
rect 12103 9356 12113 9412
rect 10496 9219 10580 9224
rect 10496 9019 10506 9219
rect 10570 9019 10580 9219
rect 10496 9014 10580 9019
rect 9026 8287 9036 8387
rect 9100 8287 9110 8387
rect 9026 8282 9110 8287
rect 10496 8388 10580 8440
rect 10496 8288 10506 8388
rect 10570 8288 10580 8388
rect 10496 8283 10580 8288
rect 8354 8275 8438 8280
rect 8354 8255 8364 8275
rect 4518 8124 4713 8129
rect 5193 8211 8364 8255
rect 8428 8211 8438 8275
rect 5193 8186 8438 8211
rect 5193 7676 5267 8186
rect 9103 8171 9283 8176
rect 9103 8107 9113 8171
rect 9273 8107 9283 8171
rect 9103 8102 9283 8107
rect 10075 8173 10255 8178
rect 10075 8109 10085 8173
rect 10245 8109 10255 8173
rect 10075 8104 10255 8109
rect 10075 7677 10139 8104
rect 8707 7676 10139 7677
rect 5193 7671 10139 7676
rect 5193 7607 5450 7671
rect 5514 7613 10139 7671
rect 5514 7607 5566 7613
rect 5193 7602 5566 7607
rect 5193 6132 5267 7602
rect 8288 7548 8438 7553
rect 8288 7484 8364 7548
rect 8428 7484 8438 7548
rect 8288 7479 8438 7484
rect 8710 6960 8784 7613
rect 5440 6955 5580 6960
rect 5440 6891 5450 6955
rect 5514 6891 5580 6955
rect 5440 6886 5580 6891
rect 8354 6955 8784 6960
rect 8354 6891 8364 6955
rect 8428 6891 8784 6955
rect 8354 6886 8784 6891
rect 8306 6239 8443 6244
rect 8306 6175 8364 6239
rect 8428 6175 8443 6239
rect 8306 6170 8443 6175
rect 5193 6127 5524 6132
rect 5193 6063 5450 6127
rect 5514 6063 5524 6127
rect 5193 6058 5524 6063
rect 5482 2402 5847 2407
rect 2985 2035 2991 2402
rect 3356 2401 5848 2402
rect 3356 2036 5482 2401
rect 5847 2036 5848 2401
rect 3356 2035 5848 2036
rect 5482 2030 5847 2035
rect 12025 1365 12113 9356
rect 13137 9412 13225 9417
rect 13137 9356 13147 9412
rect 13215 9356 13225 9412
rect 13137 8729 13225 9356
rect 13127 8634 13137 8729
rect 13225 8634 13235 8729
rect 26456 8168 26877 8173
rect 26456 7617 26466 8168
rect 26867 7617 26877 8168
rect 26456 7612 26877 7617
rect 27224 5535 27424 5540
rect 27224 5380 27234 5535
rect 27414 5380 27424 5535
rect 24729 5371 24805 5376
rect 27224 5375 27424 5380
rect 24729 5290 24739 5371
rect 24568 5206 24739 5290
rect 17855 5134 18051 5136
rect 17855 5070 17865 5134
rect 18041 5070 18051 5134
rect 17855 5068 18051 5070
rect 21643 4865 21719 4870
rect 21643 4017 21653 4865
rect 20726 3865 21653 4017
rect 21709 3865 21719 4865
rect 20726 3860 21719 3865
rect 18704 3039 18794 3044
rect 18704 2674 18714 3039
rect 17855 2669 18714 2674
rect 17855 2611 17865 2669
rect 18041 2611 18714 2669
rect 17855 2607 18714 2611
rect 18784 2607 18794 3039
rect 17855 2606 18794 2607
rect 13740 2396 16053 2401
rect 13740 2181 13750 2396
rect 16043 2181 16053 2396
rect 13740 2176 16053 2181
rect 18704 2092 18794 2606
rect 19592 3039 19683 3044
rect 19592 2607 19602 3039
rect 19673 2607 19683 3039
rect 19592 2602 19683 2607
rect 18694 2087 18804 2092
rect 18694 1988 18704 2087
rect 18794 1988 18804 2087
rect 18694 1983 18804 1988
rect 7914 1185 12113 1365
rect 7914 785 8094 1185
rect 19496 839 19697 844
rect 7904 620 7914 785
rect 8094 620 8104 785
rect 19496 690 19506 839
rect 19687 690 19697 839
rect 19496 685 19697 690
rect 20726 841 20883 3860
rect 24568 3715 24652 5206
rect 24729 5203 24739 5206
rect 24795 5203 24805 5371
rect 24729 5198 24805 5203
rect 24568 2815 24578 3715
rect 24642 2815 24652 3715
rect 24568 2810 24652 2815
rect 21013 2403 21338 2408
rect 21013 2035 21023 2403
rect 21328 2035 21338 2403
rect 21013 2030 21338 2035
rect 24333 1577 24485 1582
rect 24333 1428 24343 1577
rect 24475 1428 24485 1577
rect 24333 1423 24485 1428
rect 20726 684 23370 841
rect 23550 684 23556 841
rect 11768 678 11968 683
rect 11768 601 11778 678
rect 11958 601 11968 678
rect 15632 455 15832 460
rect 15632 385 15642 455
rect 15822 385 15832 455
<< via3 >>
rect 17732 36730 17796 42754
rect 24628 36732 24692 42756
rect 10602 30806 10666 30906
rect 2046 30057 2446 30457
rect 17731 30274 17795 36298
rect 24627 30272 24691 36296
rect 25088 29859 25439 30171
rect 11068 29599 11226 29793
rect 6236 27582 7095 27983
rect 5500 24045 5598 24115
rect 11109 21845 11209 21945
rect 22084 21556 22148 27080
rect 20127 20949 20227 21049
rect 6169 19587 6246 19687
rect 5273 19385 5373 19462
rect 19815 18439 19879 19039
rect 21403 18732 21503 18796
rect 6342 17439 6406 17639
rect 11431 17063 11495 17663
rect 11431 16035 11495 16635
rect 22084 15370 22148 20894
rect 19815 14792 19879 15259
rect 21526 14464 22053 14471
rect 21526 13980 22054 14464
rect 21526 13979 22053 13980
rect 9591 12927 10125 13059
rect 5273 11053 5373 11125
rect 6170 10327 6234 10562
rect 4365 9818 4498 9919
rect 3925 9668 4058 9768
rect 7644 9285 7708 9520
rect 9036 10104 9100 10304
rect 12349 11926 12894 12101
rect 2868 8129 3266 8529
rect 7643 8675 7709 8739
rect 5450 8323 5514 8387
rect 6161 8322 6244 8388
rect 10506 9019 10570 9219
rect 10506 8288 10570 8388
rect 9113 8107 9273 8171
rect 8364 7484 8428 7548
rect 5450 6891 5514 6955
rect 8364 6175 8428 6239
rect 2991 2035 3356 2402
rect 5482 2036 5847 2401
rect 13137 8634 13225 8729
rect 26466 7617 26867 8168
rect 27234 5380 27414 5535
rect 17865 5131 18041 5134
rect 17865 5073 18041 5131
rect 17865 5070 18041 5073
rect 13750 2181 16043 2396
rect 19602 2607 19673 3039
rect 7914 620 8094 785
rect 19506 690 19687 839
rect 21023 2035 21328 2403
rect 24343 1428 24475 1577
rect 23370 684 23550 841
rect 11778 611 11958 678
rect 11778 601 11958 611
rect 15642 395 15822 455
rect 15642 385 15822 395
<< mimcap >>
rect 11484 42702 17484 42742
rect 11484 36782 11524 42702
rect 17444 36782 17484 42702
rect 11484 36742 17484 36782
rect 18380 42704 24380 42744
rect 18380 36784 18420 42704
rect 24340 36784 24380 42704
rect 18380 36744 24380 36784
rect 11483 36246 17483 36286
rect 11483 30326 11523 36246
rect 17443 30326 17483 36246
rect 11483 30286 17483 30326
rect 18379 36244 24379 36284
rect 18379 30324 18419 36244
rect 24339 30324 24379 36244
rect 18379 30284 24379 30324
rect 22396 27028 27896 27068
rect 22396 21608 22436 27028
rect 27856 21608 27896 27028
rect 22396 21568 27896 21608
rect 22396 20842 27896 20882
rect 22396 15422 22436 20842
rect 27856 15422 27896 20842
rect 22396 15382 27896 15422
<< mimcapcontact >>
rect 11524 36782 17444 42702
rect 18420 36784 24340 42704
rect 11523 30326 17443 36246
rect 18419 30324 24339 36244
rect 22436 21608 27856 27028
rect 22436 15422 27856 20842
<< metal4 >>
rect 800 43931 1200 44152
rect 800 43741 1283 43931
rect 800 30457 1200 43741
rect 17716 42754 17812 42770
rect 11523 42702 17445 42703
rect 11523 36782 11524 42702
rect 17444 36782 17445 42702
rect 11523 36781 17445 36782
rect 16588 36247 17165 36781
rect 17716 36730 17732 42754
rect 17796 36730 17812 42754
rect 24612 42756 24708 42772
rect 18419 42704 24341 42705
rect 18419 36784 18420 42704
rect 24340 36784 24341 42704
rect 18419 36783 24341 36784
rect 17716 36714 17812 36730
rect 17715 36298 17811 36314
rect 11522 36246 17444 36247
rect 11522 30907 11523 36246
rect 10601 30906 11523 30907
rect 10601 30806 10602 30906
rect 10666 30806 11523 30906
rect 10601 30805 11523 30806
rect 2045 30457 2447 30458
rect 800 30057 2046 30457
rect 2446 30057 2447 30457
rect 800 27982 1200 30057
rect 2045 30056 2447 30057
rect 11068 29794 11226 30805
rect 11522 30326 11523 30805
rect 17443 30326 17444 36246
rect 11522 30325 17444 30326
rect 16884 29900 17437 30325
rect 17715 30274 17731 36298
rect 17795 30274 17811 36298
rect 18825 36245 19402 36783
rect 24612 36732 24628 42756
rect 24692 36732 24708 42756
rect 24612 36716 24708 36732
rect 24611 36296 24707 36312
rect 18418 36244 24340 36245
rect 18418 30324 18419 36244
rect 24339 30324 24340 36244
rect 18418 30323 24340 30324
rect 17715 30258 17811 30274
rect 18428 29900 18981 30323
rect 24611 30272 24627 36296
rect 24691 30272 24707 36296
rect 24611 30256 24707 30272
rect 25087 30171 25440 30172
rect 28400 30171 28800 44152
rect 11067 29793 11227 29794
rect 11067 29599 11068 29793
rect 11226 29599 11227 29793
rect 11067 29598 11227 29599
rect 16884 29270 18994 29900
rect 25087 29859 25088 30171
rect 25439 29859 28800 30171
rect 25087 29858 25440 29859
rect 6235 27983 7096 27984
rect 6235 27982 6236 27983
rect 800 27582 6236 27982
rect 7095 27582 7096 27983
rect 800 8529 1200 27582
rect 6235 27581 7096 27582
rect 22068 27080 22164 27096
rect 5499 24115 5599 24116
rect 4365 24045 5500 24115
rect 5598 24045 5642 24115
rect 4365 9920 4498 24045
rect 5499 24044 5599 24045
rect 11108 21945 11210 21946
rect 11108 21845 11109 21945
rect 11209 21845 11210 21945
rect 11108 21844 11210 21845
rect 6168 19687 6247 19688
rect 6008 19587 6169 19687
rect 6246 19587 6256 19687
rect 5272 19462 5374 19463
rect 5272 19385 5273 19462
rect 5373 19385 5374 19462
rect 5272 19384 5374 19385
rect 5273 11126 5373 19384
rect 6008 17640 6108 19587
rect 6168 19586 6247 19587
rect 6008 17639 6407 17640
rect 6008 17540 6342 17639
rect 6341 17439 6342 17540
rect 6406 17439 6407 17639
rect 6341 17438 6407 17439
rect 11109 17162 11209 21844
rect 22068 21556 22084 27080
rect 22148 21556 22164 27080
rect 22068 21540 22164 21556
rect 22435 27028 27857 27029
rect 22435 21608 22436 27028
rect 27856 21608 27857 27028
rect 22435 21607 27857 21608
rect 22435 21253 22936 21607
rect 21402 21151 22936 21253
rect 20126 21049 20228 21050
rect 20126 20949 20127 21049
rect 20227 20949 20228 21049
rect 20126 20948 20228 20949
rect 19814 19039 19880 19040
rect 19814 18439 19815 19039
rect 19879 18538 19880 19039
rect 20127 18538 20227 20948
rect 21402 18796 21504 21151
rect 21402 18732 21403 18796
rect 21503 18732 21504 18796
rect 21402 18731 21504 18732
rect 22068 20894 22164 20910
rect 19879 18439 20227 18538
rect 19814 18438 20227 18439
rect 11430 17663 11496 17664
rect 11430 17162 11431 17663
rect 11109 17063 11431 17162
rect 11495 17063 11496 17663
rect 11109 17062 11496 17063
rect 11109 15260 11209 17062
rect 20127 16636 20227 18438
rect 11430 16635 20227 16636
rect 11430 16035 11431 16635
rect 11495 16536 20227 16635
rect 11495 16035 11496 16536
rect 11430 16034 11496 16035
rect 22068 15370 22084 20894
rect 22148 15370 22164 20894
rect 22435 20843 22936 21151
rect 22435 20842 27857 20843
rect 22435 15422 22436 20842
rect 27856 15422 27857 20842
rect 22435 15421 27857 15422
rect 22068 15354 22164 15370
rect 11109 15259 19880 15260
rect 11109 15160 19815 15259
rect 19814 14792 19815 15160
rect 19879 14792 19880 15259
rect 19814 14782 19880 14792
rect 9591 14471 22127 14474
rect 9591 13981 21526 14471
rect 22053 14464 22127 14471
rect 28400 14464 28800 29859
rect 9591 13060 10125 13981
rect 12077 13974 12894 13981
rect 21525 13979 21526 13981
rect 22054 13981 28800 14464
rect 22054 13980 22055 13981
rect 22053 13979 22055 13980
rect 21525 13978 22054 13979
rect 9590 13059 10126 13060
rect 9590 12927 9591 13059
rect 10125 12927 10126 13059
rect 9590 12926 10126 12927
rect 12349 12102 12894 13974
rect 12348 12101 12895 12102
rect 12348 11926 12349 12101
rect 12894 11926 12895 12101
rect 12348 11925 12895 11926
rect 5272 11125 5374 11126
rect 5272 11053 5273 11125
rect 5373 11053 5374 11125
rect 5272 11052 5374 11053
rect 6169 10562 8084 10563
rect 6169 10327 6170 10562
rect 6234 10483 8084 10562
rect 6234 10327 6235 10483
rect 6169 10326 6235 10327
rect 4364 9919 4499 9920
rect 4364 9818 4365 9919
rect 4498 9818 4499 9919
rect 4364 9817 4499 9818
rect 3924 9768 4059 9769
rect 3924 9668 3925 9768
rect 4058 9668 4059 9768
rect 3924 9667 4059 9668
rect 2867 8529 3267 8530
rect 800 8129 2868 8529
rect 3266 8129 3267 8529
rect 800 2402 1200 8129
rect 2867 8128 3267 8129
rect 2990 2402 3357 2403
rect 800 2035 2991 2402
rect 3356 2035 3357 2402
rect 800 1000 1200 2035
rect 2990 2034 3357 2035
rect 3925 1561 4058 9667
rect 7984 9521 8084 10483
rect 9035 10304 9101 10305
rect 9035 10104 9036 10304
rect 9100 10167 9101 10304
rect 9100 10104 10855 10167
rect 9035 10103 10855 10104
rect 7643 9520 8084 9521
rect 7643 9285 7644 9520
rect 7708 9421 8084 9520
rect 7708 9285 7709 9421
rect 7643 8740 7709 9285
rect 10505 9219 10571 9220
rect 10505 9019 10506 9219
rect 10570 9082 10571 9219
rect 10791 9082 10855 10103
rect 10570 9019 10855 9082
rect 10505 9018 10855 9019
rect 7642 8739 7710 8740
rect 7642 8675 7643 8739
rect 7709 8675 7710 8739
rect 7642 8674 7710 8675
rect 10505 8729 10571 9018
rect 13136 8729 13226 8730
rect 10505 8634 13137 8729
rect 13225 8634 13226 8729
rect 6160 8388 6245 8389
rect 10505 8388 10571 8634
rect 13136 8633 13226 8634
rect 5449 8387 6161 8388
rect 5449 8323 5450 8387
rect 5514 8323 6161 8387
rect 5449 8322 6161 8323
rect 6244 8322 8675 8388
rect 6160 8321 6245 8322
rect 8609 7549 8675 8322
rect 10505 8288 10506 8388
rect 10570 8288 10571 8388
rect 10505 8287 10571 8288
rect 5097 7548 8675 7549
rect 5097 7484 8364 7548
rect 8428 7484 8675 7548
rect 5097 7483 8675 7484
rect 5097 6956 5163 7483
rect 5097 6955 5515 6956
rect 5097 6891 5450 6955
rect 5514 6891 5515 6955
rect 5097 6890 5515 6891
rect 8609 6864 8675 7483
rect 9112 8171 9274 8172
rect 9112 8107 9113 8171
rect 9273 8107 9274 8171
rect 9112 8106 9274 8107
rect 26465 8168 26868 8169
rect 28400 8168 28800 13981
rect 9112 6864 9176 8106
rect 26465 7617 26466 8168
rect 26867 7617 28800 8168
rect 26465 7616 26868 7617
rect 8609 6800 9176 6864
rect 8609 6240 8675 6800
rect 8362 6239 8675 6240
rect 8362 6175 8364 6239
rect 8428 6175 8675 6239
rect 8362 6174 8675 6175
rect 27233 5535 27415 5536
rect 27233 5380 27234 5535
rect 27414 5380 27415 5535
rect 27233 5379 27415 5380
rect 17864 5134 19675 5135
rect 17864 5070 17865 5134
rect 18041 5070 19675 5134
rect 17864 5069 19675 5070
rect 19599 3039 19675 5069
rect 19599 2609 19602 3039
rect 19601 2607 19602 2609
rect 19673 2609 19675 3039
rect 19673 2607 19674 2609
rect 19601 2606 19674 2607
rect 21022 2403 21329 2404
rect 21022 2402 21023 2403
rect 5481 2401 21023 2402
rect 5481 2036 5482 2401
rect 5847 2396 21023 2401
rect 5847 2181 13750 2396
rect 16043 2181 21023 2396
rect 5847 2036 21023 2181
rect 5481 2035 21023 2036
rect 21328 2402 21329 2403
rect 21328 2035 21335 2402
rect 21022 2034 21329 2035
rect 24342 1577 24476 1578
rect 24342 1561 24343 1577
rect 3925 1428 24343 1561
rect 24475 1428 24476 1577
rect 24342 1427 24476 1428
rect 24343 1418 24476 1427
rect 19506 840 19687 903
rect 23369 841 23551 842
rect 19505 839 19688 840
rect 7913 785 8095 786
rect 7913 620 7914 785
rect 8094 620 8095 785
rect 19505 690 19506 839
rect 19687 690 19688 839
rect 19505 689 19688 690
rect 7913 619 8095 620
rect 11777 678 11959 679
rect 7914 0 8094 619
rect 11777 601 11778 678
rect 11958 601 11959 678
rect 11777 600 11959 601
rect 11778 0 11958 600
rect 15641 455 15823 456
rect 15641 385 15642 455
rect 15822 385 15823 455
rect 15641 384 15823 385
rect 15642 0 15822 384
rect 19506 188 19687 689
rect 23369 684 23370 841
rect 23550 684 23551 841
rect 23369 683 23551 684
rect 19506 0 19686 188
rect 23370 0 23550 683
rect 27234 0 27414 5379
rect 28400 1000 28800 7617
<< labels >>
flabel metal4 s 27234 0 27414 200 0 FreeSans 960 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 23370 0 23550 200 0 FreeSans 960 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 19506 0 19686 200 0 FreeSans 960 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 15642 0 15822 200 0 FreeSans 960 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 11778 0 11958 200 0 FreeSans 960 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 7914 0 8094 200 0 FreeSans 960 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 800 1000 1200 44152 1 FreeSans 400 0 0 0 VGND
port 52 nsew ground bidirectional
flabel metal4 28400 1000 28800 44152 1 FreeSans 400 0 0 0 VAPWR
port 53 nsew power bidirectional
rlabel metal2 26893 5465 26893 5465 3 VCR_0.LED
rlabel metal2 26932 8128 26932 8128 3 VCR_0.vcc
rlabel metal2 21148 1871 21148 1871 7 VCR_0.Vled
rlabel metal2 24402 1555 24402 1555 5 VCR_0.VT
rlabel metal2 21114 3179 21114 3179 7 VCR_0.vss
rlabel metal3 21105 3938 21105 3938 7 VCR_0.vsen
rlabel metal2 20552 9620 20552 9620 3 Timming_0.Vd
rlabel metal2 13608 2311 13608 2311 7 Timming_0.vss
rlabel metal2 18104 2087 18104 2087 5 Timming_0.vb2
rlabel metal2 18431 2102 18431 2102 5 Timming_0.vb3
rlabel metal3 18760 2080 18760 2080 5 Timming_0.Vled
rlabel metal2 13003 11058 13003 11058 3 latch_sch_0.VDD
rlabel metal2 11231 9218 11231 9218 7 latch_sch_0.VSS
rlabel metal3 12068 9074 12068 9074 5 latch_sch_0.S
rlabel metal3 13177 9070 13177 9070 5 latch_sch_0.R
rlabel metal2 12926 10324 12926 10324 3 latch_sch_0.Q
rlabel metal2 11827 10200 11827 10200 7 latch_sch_0.Qn
rlabel metal2 10760 30190 10760 30190 5 delay_1_0.vcc
rlabel metal4 11134 29985 11134 29985 5 delay_1_0.vd_n
rlabel metal2 2325 30148 2325 30148 7 delay_1_0.vss
rlabel metal3 2819 29913 2819 29913 5 delay_1_0.vd
rlabel metal2 10812 12779 10812 12779 3 COMP_2_0.vcc
rlabel metal2 5273 5769 5273 5769 7 COMP_2_0.vss
rlabel metal2 5668 9712 5668 9712 7 COMP_2_0.vin_p
rlabel metal4 10900 8681 10900 8681 3 COMP_2_0.out
rlabel metal2 5668 9869 5668 9869 1 COMP_2_0.vin_n
rlabel metal2 5726 11089 5726 11089 7 COMP_2_0.vb
rlabel metal2 7735 12058 7735 12058 7 COMP_2_0.vd_n
rlabel metal2 7962 14074 7962 14074 7 BIAS_1_0.vcc
rlabel metal1 17792 28262 17792 28262 3 BIAS_1_0.vss
rlabel metal2 7988 14913 7988 14913 7 BIAS_1_0.vd_n
rlabel metal2 5938 19435 5938 19435 7 BIAS_1_0.vb
rlabel metal3 5663 24075 5663 24075 7 BIAS_1_0.vth
flabel locali 16847 27558 17095 27662 0 FreeSans 400 0 0 0 BIAS_1_0.XQ12.Emitter
flabel locali 16935 26987 17036 27036 0 FreeSans 400 0 0 0 BIAS_1_0.XQ12.Collector
flabel locali 16941 27146 17059 27186 0 FreeSans 400 0 0 0 BIAS_1_0.XQ12.Base
flabel locali 16847 26214 17095 26318 0 FreeSans 400 0 0 0 BIAS_1_0.XQ11.Emitter
flabel locali 16935 25643 17036 25692 0 FreeSans 400 0 0 0 BIAS_1_0.XQ11.Collector
flabel locali 16941 25802 17059 25842 0 FreeSans 400 0 0 0 BIAS_1_0.XQ11.Base
flabel locali 14159 27558 14407 27662 0 FreeSans 400 0 0 0 BIAS_1_0.XQ10.Emitter
flabel locali 14247 26987 14348 27036 0 FreeSans 400 0 0 0 BIAS_1_0.XQ10.Collector
flabel locali 14253 27146 14371 27186 0 FreeSans 400 0 0 0 BIAS_1_0.XQ10.Base
flabel locali 15503 27558 15751 27662 0 FreeSans 400 0 0 0 BIAS_1_0.XQ9.Emitter
flabel locali 15591 26987 15692 27036 0 FreeSans 400 0 0 0 BIAS_1_0.XQ9.Collector
flabel locali 15597 27146 15715 27186 0 FreeSans 400 0 0 0 BIAS_1_0.XQ9.Base
flabel locali 14159 26214 14407 26318 0 FreeSans 400 0 0 0 BIAS_1_0.XQ8.Emitter
flabel locali 14247 25643 14348 25692 0 FreeSans 400 0 0 0 BIAS_1_0.XQ8.Collector
flabel locali 14253 25802 14371 25842 0 FreeSans 400 0 0 0 BIAS_1_0.XQ8.Base
flabel locali 16847 24870 17095 24974 0 FreeSans 400 0 0 0 BIAS_1_0.XQ7.Emitter
flabel locali 16935 24299 17036 24348 0 FreeSans 400 0 0 0 BIAS_1_0.XQ7.Collector
flabel locali 16941 24458 17059 24498 0 FreeSans 400 0 0 0 BIAS_1_0.XQ7.Base
flabel locali 14159 24870 14407 24974 0 FreeSans 400 0 0 0 BIAS_1_0.XQ6.Emitter
flabel locali 14247 24299 14348 24348 0 FreeSans 400 0 0 0 BIAS_1_0.XQ6.Collector
flabel locali 14253 24458 14371 24498 0 FreeSans 400 0 0 0 BIAS_1_0.XQ6.Base
flabel locali 15503 24870 15751 24974 0 FreeSans 400 0 0 0 BIAS_1_0.XQ5.Emitter
flabel locali 15591 24299 15692 24348 0 FreeSans 400 0 0 0 BIAS_1_0.XQ5.Collector
flabel locali 15597 24458 15715 24498 0 FreeSans 400 0 0 0 BIAS_1_0.XQ5.Base
flabel locali 15503 26214 15751 26318 0 FreeSans 400 0 0 0 BIAS_1_0.XQ4.Emitter
flabel locali 15591 25643 15692 25692 0 FreeSans 400 0 0 0 BIAS_1_0.XQ4.Collector
flabel locali 15597 25802 15715 25842 0 FreeSans 400 0 0 0 BIAS_1_0.XQ4.Base
<< end >>
